module DenseWeightLut #(parameter
    WORD_SIZE = 32, 
    LENGTH_SIZE = 10,
    ADR_SIZE = 4
) (
    clk,
    adr,
    dataOut
);

    input                   clk;
    input   [ADR_SIZE-1:0]  adr;
    output  [WORD_SIZE-1:0] dataOut;

    wire [WORD_SIZE-1:0] mem [0:LENGTH_SIZE-1];

    assign dataOut = mem[adr];

    assign mem[0] = 32'b11110011001111111111011101000000;
   assign mem[1] = 32'b11111010000001101111101000101000;
   assign mem[2] = 32'b00000010001111010010011101111100;
   assign mem[3] = 32'b00001101010100001111111011110000;
   assign mem[4] = 32'b00000111010101011001101000010000;
   assign mem[5] = 32'b11110100011101011101011011000000;
   assign mem[6] = 32'b00000010001001101100110010101000;
   assign mem[7] = 32'b00000101011110010111100011000000;
   assign mem[8] = 32'b11111000011111110001101011000000;
   assign mem[9] = 32'b11110001010101100110110000110000;
   assign mem[10] = 32'b11111010101110111000000010011000;
   assign mem[11] = 32'b00000000011011110110101110100010;
   assign mem[12] = 32'b00010000001101101011110110100000;
   assign mem[13] = 32'b11111000001111011111110110111000;
   assign mem[14] = 32'b00000010011011000111011010100000;
   assign mem[15] = 32'b11111111000000001111011001101000;
   assign mem[16] = 32'b00001011111001010000000101110000;
   assign mem[17] = 32'b11111101011011110010010100111000;
   assign mem[18] = 32'b11110010110000110000011001010000;
   assign mem[19] = 32'b11110110110000010100110111010000;
   assign mem[20] = 32'b11111101011100101110001011010000;
   assign mem[21] = 32'b00001010110000001000110001010000;
   assign mem[22] = 32'b11110110011000001111010001110000;
   assign mem[23] = 32'b00000101100000101010011111100000;
   assign mem[24] = 32'b00000111011101001000101101010000;
   assign mem[25] = 32'b11111110110001110000000111000100;
   assign mem[26] = 32'b00000000110001110101001110001100;
   assign mem[27] = 32'b00000000101010010101010001000100;
   assign mem[28] = 32'b11111110000000111001110001001010;
   assign mem[29] = 32'b11110101101011000100110111100000;
   assign mem[30] = 32'b00000010011110101111011110111100;
   assign mem[31] = 32'b00000011111001100010001001000100;
   assign mem[32] = 32'b00001000111100011101110000110000;
   assign mem[33] = 32'b00000100001001100100010011001000;
   assign mem[34] = 32'b11111010101101011101101111010000;
   assign mem[35] = 32'b11111000010101010011001110101000;
   assign mem[36] = 32'b11111001100001100111111001000000;
   assign mem[37] = 32'b11111000010001100001001101111000;
   assign mem[38] = 32'b11110110010011110110100000110000;
   assign mem[39] = 32'b11111001100101100010011111101000;
   assign mem[40] = 32'b00000001010100111100111010000000;
   assign mem[41] = 32'b00000001100010110001111110011100;
   assign mem[42] = 32'b11111011000000011001000011000000;
   assign mem[43] = 32'b00000011000000001010010011000000;
   assign mem[44] = 32'b11111101001011111101011110110100;
   assign mem[45] = 32'b11111001001111010110100100110000;
   assign mem[46] = 32'b11111010110100001110001001110000;
   assign mem[47] = 32'b11111011110001101011101100101000;
   assign mem[48] = 32'b00000011000001110110101101100100;
   assign mem[49] = 32'b00000001100000000011111101000110;
   assign mem[50] = 32'b11111000110100011111010101100000;
   assign mem[51] = 32'b11111110001110011111001101100000;
   assign mem[52] = 32'b11110111011001010111100011110000;
   assign mem[53] = 32'b00000001010110101100111100110110;
   assign mem[54] = 32'b11111001011000100110101100110000;
   assign mem[55] = 32'b11111110100011011111011111001000;
   assign mem[56] = 32'b00000000011010011110111110110101;
   assign mem[57] = 32'b00000011100100001010101011011100;
   assign mem[58] = 32'b00001001111100101001001010010000;
   assign mem[59] = 32'b11111001111100110011011010010000;
   assign mem[60] = 32'b00000000100010111010110100110000;
   assign mem[61] = 32'b11111111001001000010110110000111;
   assign mem[62] = 32'b11111110101110001101100101010100;
   assign mem[63] = 32'b11111100101011000110100110111000;
   assign mem[64] = 32'b00000011001000110101000101000000;
   assign mem[65] = 32'b00000101010000010111010111011000;
   assign mem[66] = 32'b00000011001101001101101101010100;
   assign mem[67] = 32'b00000011011000111001000110100000;
   assign mem[68] = 32'b00000101001101111010101100000000;
   assign mem[69] = 32'b11111011111101110101001100101000;
   assign mem[70] = 32'b11111111111010111001001010100000;
   assign mem[71] = 32'b11111001101100101000001000110000;
   assign mem[72] = 32'b11111110111011111110011011011000;
   assign mem[73] = 32'b00000011111011111101111101000100;
   assign mem[74] = 32'b11111100111011111010101000000000;
   assign mem[75] = 32'b00000010001100101011110010000100;
   assign mem[76] = 32'b00000011111000101011110100000100;
   assign mem[77] = 32'b11111011101000101111111111111000;
   assign mem[78] = 32'b11110110110010100110110010100000;
   assign mem[79] = 32'b11111010111010010101011010001000;
   assign mem[80] = 32'b00000011110110000001011010110100;
   assign mem[81] = 32'b00001001000010111011010000010000;
   assign mem[82] = 32'b11111100110110010100011011000000;
   assign mem[83] = 32'b00000001101101011000001111110010;
   assign mem[84] = 32'b00000011111011111111010100010000;
   assign mem[85] = 32'b11111101100001010100000111010000;
   assign mem[86] = 32'b11111001001100000001100101100000;
   assign mem[87] = 32'b00000110001100010011010101001000;
   assign mem[88] = 32'b00000001111000011101001110101010;
   assign mem[89] = 32'b00000001011110100011111011011100;
   assign mem[90] = 32'b00000001010111100010110011000000;
   assign mem[91] = 32'b11111001101011100010111000000000;
   assign mem[92] = 32'b11111101110000110101010011010000;
   assign mem[93] = 32'b11111010001000001110110010100000;
   assign mem[94] = 32'b11111100110111101011100010010000;
   assign mem[95] = 32'b11111100000010000010111001011100;
   assign mem[96] = 32'b00000111101000100111100000110000;
   assign mem[97] = 32'b11111110100011000010110100000100;
   assign mem[98] = 32'b00000001000001111011100101111110;
   assign mem[99] = 32'b00000000101010110011110111000010;
   assign mem[100] = 32'b11111111101011111011001110011101;
   assign mem[101] = 32'b11111100011101101011011000000000;
   assign mem[102] = 32'b00000101101100000100010011110000;
   assign mem[103] = 32'b00000011111100010111110111011000;
   assign mem[104] = 32'b11111001101101110110001110010000;
   assign mem[105] = 32'b11111011101000111001111010101000;
   assign mem[106] = 32'b00001000110100111001100011100000;
   assign mem[107] = 32'b11111100110010001000011000111100;
   assign mem[108] = 32'b11111101001001001111101101111000;
   assign mem[109] = 32'b11111110011111000100111011101110;
   assign mem[110] = 32'b11110110100011011000101100110000;
   assign mem[111] = 32'b00000010101011100010100010110100;
   assign mem[112] = 32'b11111100000010100110100100101000;
   assign mem[113] = 32'b00000100100110001010010101001000;
   assign mem[114] = 32'b00000010111111001011101111100100;
   assign mem[115] = 32'b00000001010111101011000101010000;
   assign mem[116] = 32'b11111110111101111110001100000000;
   assign mem[117] = 32'b00000111101111101100011001000000;
   assign mem[118] = 32'b11111100000100100011110110100000;
   assign mem[119] = 32'b11110100001011011101110100110000;
   assign mem[120] = 32'b11111111000100001111010010001111;
   assign mem[121] = 32'b11111010010101110001001101011000;
   assign mem[122] = 32'b00000001010000100110111110011100;
   assign mem[123] = 32'b00000100001010101011000111100000;
   assign mem[124] = 32'b11111101000101000100101011111100;
   assign mem[125] = 32'b11111101000000011110011000011000;
   assign mem[126] = 32'b11110101101100110010000101100000;
   assign mem[127] = 32'b00000100010000110000001001110000;
   assign mem[128] = 32'b11111100001001111111111010111000;
   assign mem[129] = 32'b11111100111100011000000100100100;
   assign mem[130] = 32'b00000011100111110001010111011000;
   assign mem[131] = 32'b00001100110100010101100110110000;
   assign mem[132] = 32'b11110111111000111101011010110000;
   assign mem[133] = 32'b00000011000100010001110001100100;
   assign mem[134] = 32'b11111111111111010101000000000001;
   assign mem[135] = 32'b11111011000011101000001001010000;
   assign mem[136] = 32'b11110001111100110100100001010000;
   assign mem[137] = 32'b00000100000111111111011100111000;
   assign mem[138] = 32'b11111111110001011101110010101100;
   assign mem[139] = 32'b00000001110011010110000111101000;
   assign mem[140] = 32'b00000001000001010110101010111110;
   assign mem[141] = 32'b11111110110001001001111000001000;
   assign mem[142] = 32'b00000000100000010001101010011100;
   assign mem[143] = 32'b00000110110101101100101000010000;
   assign mem[144] = 32'b00000110010111000101101011101000;
   assign mem[145] = 32'b11110111010110011100111100110000;
   assign mem[146] = 32'b11111011111010011101000001001000;
   assign mem[147] = 32'b00000000110011101110000101001010;
   assign mem[148] = 32'b11111110110100011000000001111010;
   assign mem[149] = 32'b11111001111100011011110001011000;
   assign mem[150] = 32'b00000010100000100000001011100100;
   assign mem[151] = 32'b11111011000101001100011100110000;
   assign mem[152] = 32'b00000000101011011100110101011011;
   assign mem[153] = 32'b00000010001001100001110111011100;
   assign mem[154] = 32'b11111011011100000011100000010000;
   assign mem[155] = 32'b11111100100100100010010101111000;
   assign mem[156] = 32'b00000101111100001100010110111000;
   assign mem[157] = 32'b11110111111111011011110010100000;
   assign mem[158] = 32'b00000101000010110001111100010000;
   assign mem[159] = 32'b00000001111110111011101111111100;
   assign mem[160] = 32'b11110111001011111100101010000000;
   assign mem[161] = 32'b00000001010100011010110001011010;
   assign mem[162] = 32'b00001011011100010111100101000000;
   assign mem[163] = 32'b00000010010111101110011101101000;
   assign mem[164] = 32'b11111011101111010101100100111000;
   assign mem[165] = 32'b11101011010011001001111001100000;
   assign mem[166] = 32'b00000010110100100011111110000100;
   assign mem[167] = 32'b00000100011000011010111001001000;
   assign mem[168] = 32'b11110100111101010010110101110000;
   assign mem[169] = 32'b11110011010000111100001011100000;
   assign mem[170] = 32'b11111110101110011111101101000100;
   assign mem[171] = 32'b00000111100000001101100010011000;
   assign mem[172] = 32'b11111001001010001111111101001000;
   assign mem[173] = 32'b00000101011111110010011011010000;
   assign mem[174] = 32'b00000000100001010111001110100111;
   assign mem[175] = 32'b11111111011111110010110111000111;
   assign mem[176] = 32'b00000010010100100110101001011000;
   assign mem[177] = 32'b11111101100000011000010011011100;
   assign mem[178] = 32'b11111111101011100010001100011011;
   assign mem[179] = 32'b11110101001011101011111010010000;
   assign mem[180] = 32'b11111011010111011001010011001000;
   assign mem[181] = 32'b00000011100000000100100100101000;
   assign mem[182] = 32'b11111101110001100001101111110100;
   assign mem[183] = 32'b11111001101110000001000011101000;
   assign mem[184] = 32'b00001110100111100110110010010000;
   assign mem[185] = 32'b11110111100000000011011111100000;
   assign mem[186] = 32'b00000011111111010011110000100100;
   assign mem[187] = 32'b00000101001000011100010011110000;
   assign mem[188] = 32'b11101101101010101111001110100000;
   assign mem[189] = 32'b11101000011011001000110100000000;
   assign mem[190] = 32'b11111001011100100010111001111000;
   assign mem[191] = 32'b11111110000111010000111100001110;
   assign mem[192] = 32'b11111111011011011001110111000111;
   assign mem[193] = 32'b00000101000010001110100101111000;
   assign mem[194] = 32'b00001000100000011001011010110000;
   assign mem[195] = 32'b11111000110111010100111111000000;
   assign mem[196] = 32'b00000000111011011111110100011110;
   assign mem[197] = 32'b11110101100111110110010100110000;
   assign mem[198] = 32'b00000110011100000001011111001000;
   assign mem[199] = 32'b11111111010110110010010110000111;
   assign mem[200] = 32'b00000011001011110000110101101100;
   assign mem[201] = 32'b11111010100010101101101111101000;
   assign mem[202] = 32'b11111001111101110101011000110000;
   assign mem[203] = 32'b00000001010110001111110011111010;
   assign mem[204] = 32'b11111110110001011011010010001000;
   assign mem[205] = 32'b00000000000010101000011010000111;
   assign mem[206] = 32'b00001110010010101011000111010000;
   assign mem[207] = 32'b11110111101110010111101001100000;
   assign mem[208] = 32'b11111111110101100101110001010101;
   assign mem[209] = 32'b00000000111001111000000000111011;
   assign mem[210] = 32'b00000100001111001010000110001000;
   assign mem[211] = 32'b11111110101101111100010000010110;
   assign mem[212] = 32'b11111100111110000111011000101100;
   assign mem[213] = 32'b00000100110011000100000110110000;
   assign mem[214] = 32'b00000001110011001001011111011010;
   assign mem[215] = 32'b11110110011101100100011010100000;
   assign mem[216] = 32'b11111111101110001111100011010110;
   assign mem[217] = 32'b00000001100011100100111010010000;
   assign mem[218] = 32'b00000000110110101010010101011111;
   assign mem[219] = 32'b00000001111101010000101011111000;
   assign mem[220] = 32'b11110101110000111101000101010000;
   assign mem[221] = 32'b11111101110101000001100001101000;
   assign mem[222] = 32'b11111010001010101100111111000000;
   assign mem[223] = 32'b00000101010001100001001100101000;
   assign mem[224] = 32'b11111111100110100011110100010011;
   assign mem[225] = 32'b11111100001111101100100001011000;
   assign mem[226] = 32'b00001100001100101111011001110000;
   assign mem[227] = 32'b11110111000001100001110110100000;
   assign mem[228] = 32'b00000000100100101100011101000101;
   assign mem[229] = 32'b11110101101100010010110011100000;
   assign mem[230] = 32'b11111111000101000100010101111100;
   assign mem[231] = 32'b00001011100000110110111011100000;
   assign mem[232] = 32'b11110101111011100001001011100000;
   assign mem[233] = 32'b00000011001101010111100100010100;
   assign mem[234] = 32'b11111111100011011001101101100100;
   assign mem[235] = 32'b00000001011101110001000111111010;
   assign mem[236] = 32'b00001000101001000101010100010000;
   assign mem[237] = 32'b00000101000001010000101001111000;
   assign mem[238] = 32'b00000000000100001100111101111001;
   assign mem[239] = 32'b11110110101011100110010000010000;
   assign mem[240] = 32'b11111011000001011101100001000000;
   assign mem[241] = 32'b00001000111101100101000011110000;
   assign mem[242] = 32'b11110011000010010111101001000000;
   assign mem[243] = 32'b00000101010010000101111111011000;
   assign mem[244] = 32'b00000010100010110011110100111100;
   assign mem[245] = 32'b00000111001010000111101001011000;
   assign mem[246] = 32'b00000101111001100111011100101000;
   assign mem[247] = 32'b00000010110010110101111101000000;
   assign mem[248] = 32'b11111001011101010110101011100000;
   assign mem[249] = 32'b11110010111101010100110010010000;
   assign mem[250] = 32'b11111010011110010100101100000000;
   assign mem[251] = 32'b11111011101000111101010111101000;
   assign mem[252] = 32'b11111100001001111011000110011100;
   assign mem[253] = 32'b11111110101011010001010011001100;
   assign mem[254] = 32'b11111101001001100101001000001100;
   assign mem[255] = 32'b00000000101110100110111110010111;
   assign mem[256] = 32'b00001011110000111110000011110000;
   assign mem[257] = 32'b00000001100101100110001000010000;
   assign mem[258] = 32'b11111111001011011000110110011110;
   assign mem[259] = 32'b11111110101110100111101100011100;
   assign mem[260] = 32'b11101111011101111010101010100000;
   assign mem[261] = 32'b00000000110100110110100111111110;
   assign mem[262] = 32'b11111110101011111100011001111000;
   assign mem[263] = 32'b11110011001110100110110111110000;
   assign mem[264] = 32'b00000010101001001001010111011000;
   assign mem[265] = 32'b00000010000011110110011011101100;
   assign mem[266] = 32'b00001110010100111011111010010000;
   assign mem[267] = 32'b11110101100000101101010011010000;
   assign mem[268] = 32'b11111111001100110101011001100001;
   assign mem[269] = 32'b11101111111111010110010100000000;
   assign mem[270] = 32'b00000000101110001100011010101101;
   assign mem[271] = 32'b11111100101001110111000000010100;
   assign mem[272] = 32'b11111111110000110101000001011101;
   assign mem[273] = 32'b00000010100100001011010000010000;
   assign mem[274] = 32'b00000010101110011011110000100100;
   assign mem[275] = 32'b11111110010100010100111111110100;
   assign mem[276] = 32'b11111101000001001000011011111100;
   assign mem[277] = 32'b11111111001110011000101001011011;
   assign mem[278] = 32'b00000100110000100010111011000000;
   assign mem[279] = 32'b00000000100111010100101011100111;
   assign mem[280] = 32'b11111111110011001011101100000001;
   assign mem[281] = 32'b11111011100100001111100000111000;
   assign mem[282] = 32'b00000100110111001010111100001000;
   assign mem[283] = 32'b00001000100110100100100110110000;
   assign mem[284] = 32'b11111110111100010010000001000000;
   assign mem[285] = 32'b11111110101110100101001011010010;
   assign mem[286] = 32'b00000001100001110001010000101000;
   assign mem[287] = 32'b11111011011010100100110101100000;
   assign mem[288] = 32'b11111110001110010101110000101100;
   assign mem[289] = 32'b11111101001111000000111001010100;
   assign mem[290] = 32'b00000001011011010010001101110110;
   assign mem[291] = 32'b00000101011010110010001110110000;
   assign mem[292] = 32'b11111110111100011110101001001000;
   assign mem[293] = 32'b00000001100001101011010011111000;
   assign mem[294] = 32'b00000000011100001010011111110110;
   assign mem[295] = 32'b11111010001100110101011001011000;
   assign mem[296] = 32'b11111010100110001000000111110000;
   assign mem[297] = 32'b00000010001110001010100011010100;
   assign mem[298] = 32'b11111111110110110100010001100001;
   assign mem[299] = 32'b11111110110010011110010001010000;
   assign mem[300] = 32'b00000001000111110010100101111110;
   assign mem[301] = 32'b00000001011011011110010010101000;
   assign mem[302] = 32'b11111101101110111010110001001000;
   assign mem[303] = 32'b11110111001100010010111111010000;
   assign mem[304] = 32'b11111111110000111011000001110000;
   assign mem[305] = 32'b11111111011011100001011001111100;
   assign mem[306] = 32'b00001101011110100000101111110000;
   assign mem[307] = 32'b00000001001011011000000111010010;
   assign mem[308] = 32'b11111010100111010111001101100000;
   assign mem[309] = 32'b11101000100001100110000000100000;
   assign mem[310] = 32'b11111011110001011111011000101000;
   assign mem[311] = 32'b11111101010011110111000010111000;
   assign mem[312] = 32'b00000010000001110001110100100000;
   assign mem[313] = 32'b00000101100100011100100000111000;
   assign mem[314] = 32'b11111010110001000001001011100000;
   assign mem[315] = 32'b11101010101101010101101000100000;
   assign mem[316] = 32'b00000100101010011010111111101000;
   assign mem[317] = 32'b00000101011001100100100000111000;
   assign mem[318] = 32'b11110011000110000000100100100000;
   assign mem[319] = 32'b11110010111011001010111101000000;
   assign mem[320] = 32'b00000110001000101011000111011000;
   assign mem[321] = 32'b11110011001110001100000100110000;
   assign mem[322] = 32'b00000001010100011111101100101100;
   assign mem[323] = 32'b00000010000010000110100000010000;
   assign mem[324] = 32'b00000010010011101011010110100000;
   assign mem[325] = 32'b11111011111101011100111000110000;
   assign mem[326] = 32'b00000100001101001100110001101000;
   assign mem[327] = 32'b11111101011010100111010001100000;
   assign mem[328] = 32'b00000111001010101000011100100000;
   assign mem[329] = 32'b11110111011111111000001111000000;
   assign mem[330] = 32'b11111101010000000101100011001100;
   assign mem[331] = 32'b11111101010110000101010001001100;
   assign mem[332] = 32'b11111111111011000000010101110100;
   assign mem[333] = 32'b00000100010000110001011111100000;
   assign mem[334] = 32'b00000110000000001001100101001000;
   assign mem[335] = 32'b11111100100101111100110110101100;
   assign mem[336] = 32'b00001001110101001100101101100000;
   assign mem[337] = 32'b11110100000000001100010100110000;
   assign mem[338] = 32'b00000001101101000000110100100110;
   assign mem[339] = 32'b11111001111011010000010101111000;
   assign mem[340] = 32'b11110111100001100100000000110000;
   assign mem[341] = 32'b11111100000000001111010110101100;
   assign mem[342] = 32'b00000001011000001010001011111010;
   assign mem[343] = 32'b00000011011000110000101001001100;
   assign mem[344] = 32'b11111110110111110011010110010100;
   assign mem[345] = 32'b11110100110010001111111111110000;
   assign mem[346] = 32'b00001010110100111100101001000000;
   assign mem[347] = 32'b00000000111101010011010111001110;
   assign mem[348] = 32'b11110110100000000001001100010000;
   assign mem[349] = 32'b11101110001001110001001111000000;
   assign mem[350] = 32'b00000100001111101001011111100000;
   assign mem[351] = 32'b11110111101100101011111110100000;
   assign mem[352] = 32'b11111110101000101011001110101100;
   assign mem[353] = 32'b11111101110100110111000000100100;
   assign mem[354] = 32'b11111101111001100000110010100100;
   assign mem[355] = 32'b00000000001100101111000001001010;
   assign mem[356] = 32'b11111001110111100111011100101000;
   assign mem[357] = 32'b00000000000010010110011010110011;
   assign mem[358] = 32'b00001001010010110100111000010000;
   assign mem[359] = 32'b00000010101010011010110011111000;
   assign mem[360] = 32'b00000000011000100101010101101101;
   assign mem[361] = 32'b00000110111011010010101011110000;
   assign mem[362] = 32'b11111111110111110111111101101101;
   assign mem[363] = 32'b11111011010101010110110111110000;
   assign mem[364] = 32'b00000010111000011110110100101100;
   assign mem[365] = 32'b11111111111000011110000110001100;
   assign mem[366] = 32'b11110110111101101110100100100000;
   assign mem[367] = 32'b00000100011000101110100101000000;
   assign mem[368] = 32'b11111101110111010111000001100100;
   assign mem[369] = 32'b11111100111001100101110000011100;
   assign mem[370] = 32'b11111010000110011011110110111000;
   assign mem[371] = 32'b00001100010111101100101111000000;
   assign mem[372] = 32'b11110111100101000010000110010000;
   assign mem[373] = 32'b00001001000000010111101010000000;
   assign mem[374] = 32'b00000001001010101101010110011100;
   assign mem[375] = 32'b11111101111010100001100010101000;
   assign mem[376] = 32'b00000011011001110100001111101100;
   assign mem[377] = 32'b00001010011001000011001001100000;
   assign mem[378] = 32'b11111110011001000001111011100110;
   assign mem[379] = 32'b11110101000110101101001111010000;
   assign mem[380] = 32'b00000001011011111110111110100000;
   assign mem[381] = 32'b11111111111001010011010111000000;
   assign mem[382] = 32'b00000000100000011000111100011100;
   assign mem[383] = 32'b00000111011111110110101111010000;
   assign mem[384] = 32'b11111010000110111010001101110000;
   assign mem[385] = 32'b11111011000000111110101001000000;
   assign mem[386] = 32'b00000000110101101000110000101110;
   assign mem[387] = 32'b00000101111111011110101001111000;
   assign mem[388] = 32'b11110111011101100001010111100000;
   assign mem[389] = 32'b11111110111110101110101010011100;
   assign mem[390] = 32'b00000111001011100101110010111000;
   assign mem[391] = 32'b11111010010110111010001111001000;
   assign mem[392] = 32'b11111101011010110010101000111000;
   assign mem[393] = 32'b00000000100110100011001011000110;
   assign mem[394] = 32'b11111100101011110010010010101100;
   assign mem[395] = 32'b11111110100111100111011101011010;
   assign mem[396] = 32'b11111000000001001111110001010000;
   assign mem[397] = 32'b11111100110010110000001110010100;
   assign mem[398] = 32'b11111101000100100010001110011000;
   assign mem[399] = 32'b00000001111110111110011110101000;
   assign mem[400] = 32'b11111100011111001010001100010000;
   assign mem[401] = 32'b00001001110011010111101101010000;
   assign mem[402] = 32'b11111100011001001001101110101100;
   assign mem[403] = 32'b00000001111001000000001011011100;
   assign mem[404] = 32'b00000011110001110100110111000100;
   assign mem[405] = 32'b11111000011110101000110010111000;
   assign mem[406] = 32'b11111001000111111001000001110000;
   assign mem[407] = 32'b11111110110110000011110011010100;
   assign mem[408] = 32'b11111010110010000111100100011000;
   assign mem[409] = 32'b11110101000101100100011101010000;
   assign mem[410] = 32'b11110110111000001000111001110000;
   assign mem[411] = 32'b11111100001000110110100011110100;
   assign mem[412] = 32'b00000010110111001110000011101000;
   assign mem[413] = 32'b00000101011101001001010010111000;
   assign mem[414] = 32'b11110111110011011111101100100000;
   assign mem[415] = 32'b11110010000010100011001110100000;
   assign mem[416] = 32'b11111011000000110001110011001000;
   assign mem[417] = 32'b11111001001011111000010101010000;
   assign mem[418] = 32'b11111001010100111011101001100000;
   assign mem[419] = 32'b00000000111010100001011110111011;
   assign mem[420] = 32'b11111001111100010100110101011000;
   assign mem[421] = 32'b00000011010101001011100101000100;
   assign mem[422] = 32'b00000001100111101010001110000110;
   assign mem[423] = 32'b00000101100110110000101010010000;
   assign mem[424] = 32'b11111101100010011010000101010000;
   assign mem[425] = 32'b11101111001010010001010101100000;
   assign mem[426] = 32'b00000010010100110000101011011100;
   assign mem[427] = 32'b00000101010000011000101000000000;
   assign mem[428] = 32'b00000010110110111000011100010100;
   assign mem[429] = 32'b11111100100110010001010100100000;
   assign mem[430] = 32'b11110100111100110010101011110000;
   assign mem[431] = 32'b00000001100100001010011100111110;
   assign mem[432] = 32'b00000000101011101110110111111000;
   assign mem[433] = 32'b11111001101001110110001000100000;
   assign mem[434] = 32'b11111110101011101001111011011010;
   assign mem[435] = 32'b11111110011010010101011111101000;
   assign mem[436] = 32'b00010001100001011001101001000000;
   assign mem[437] = 32'b11111101010000000000110000010000;
   assign mem[438] = 32'b11111110001000010001100100011000;
   assign mem[439] = 32'b11111110010111100001100100101000;
   assign mem[440] = 32'b00000001000000111000000001110100;
   assign mem[441] = 32'b00000011010100000100011001010000;
   assign mem[442] = 32'b11111111101000001101110110000000;
   assign mem[443] = 32'b00000110010100010000101000011000;
   assign mem[444] = 32'b11111000010100000001110010011000;
   assign mem[445] = 32'b11111010000100000100101110111000;
   assign mem[446] = 32'b11111110011001110110111010001000;
   assign mem[447] = 32'b00000000101110010011111101001011;
   assign mem[448] = 32'b11111100101100000010100111000100;
   assign mem[449] = 32'b11111101101101101000111011000100;
   assign mem[450] = 32'b00000100010011011010000001101000;
   assign mem[451] = 32'b11111100100100010100111011111000;
   assign mem[452] = 32'b11111100011000010110000101001100;
   assign mem[453] = 32'b11111111100110000010001110011010;
   assign mem[454] = 32'b00000100010000000100001001101000;
   assign mem[455] = 32'b11111111111011111100000100100100;
   assign mem[456] = 32'b00000001000100010010110111101110;
   assign mem[457] = 32'b00000101101100001110010011001000;
   assign mem[458] = 32'b11111111101000101011000110111110;
   assign mem[459] = 32'b11111011011011001110001011011000;
   assign mem[460] = 32'b11111110000100010100001011110000;
   assign mem[461] = 32'b11110100001110100011100101000000;
   assign mem[462] = 32'b00000001100000001110001100100110;
   assign mem[463] = 32'b11111000010111110010010010110000;
   assign mem[464] = 32'b11111111110101111110010101110111;
   assign mem[465] = 32'b00000011101010001011111101111000;
   assign mem[466] = 32'b00001011110000010000111000010000;
   assign mem[467] = 32'b11111100011110111100011001010100;
   assign mem[468] = 32'b00000000110011111000100100110111;
   assign mem[469] = 32'b00000000011001011011010000101101;
   assign mem[470] = 32'b00000000100101011101010111010011;
   assign mem[471] = 32'b00000000111100011101011000001000;
   assign mem[472] = 32'b00000001101100000011011111110110;
   assign mem[473] = 32'b11111101101111001011010111000000;
   assign mem[474] = 32'b11111100111100101010111101011000;
   assign mem[475] = 32'b11111011101111101001111110111000;
   assign mem[476] = 32'b00000010100111010011010011111100;
   assign mem[477] = 32'b11111101110000000010101000000100;
   assign mem[478] = 32'b11111111101011010101010100000100;
   assign mem[479] = 32'b11111100111110110010000101011100;
   assign mem[480] = 32'b11111100110111000011101100110000;
   assign mem[481] = 32'b11111100010111110100000000010000;
   assign mem[482] = 32'b00000001110101000111100100111010;
   assign mem[483] = 32'b00000100010110100110110001010000;
   assign mem[484] = 32'b11111110000101010111100101101100;
   assign mem[485] = 32'b11111010111110011000110111000000;
   assign mem[486] = 32'b00000001011111000100101001010110;
   assign mem[487] = 32'b11111110110101100011110100111100;
   assign mem[488] = 32'b11111011011101111000011111000000;
   assign mem[489] = 32'b11111101111001100100100011001100;
   assign mem[490] = 32'b00000000001000011000111001100101;
   assign mem[491] = 32'b11110111110010011111001111110000;
   assign mem[492] = 32'b11111111000110111010011001000100;
   assign mem[493] = 32'b00000011001011011001101110100100;
   assign mem[494] = 32'b11111011011010001111100101100000;
   assign mem[495] = 32'b11111111100100101111101001011010;
   assign mem[496] = 32'b00001000100001001010001101110000;
   assign mem[497] = 32'b11111010100010010101001101011000;
   assign mem[498] = 32'b00000101110011010101000000000000;
   assign mem[499] = 32'b11111010010100000111000100110000;
   assign mem[500] = 32'b11111010001001011010100100001000;
   assign mem[501] = 32'b11111000110000101101101100010000;
   assign mem[502] = 32'b00000011010100100001111010111000;
   assign mem[503] = 32'b00000110010001100111010011010000;
   assign mem[504] = 32'b00001001000000001001101101110000;
   assign mem[505] = 32'b11111010010000100101100011010000;
   assign mem[506] = 32'b00000010101000111100110001110000;
   assign mem[507] = 32'b11101111001100001011100100100000;
   assign mem[508] = 32'b00000010110000001111101001011000;
   assign mem[509] = 32'b00000000010101011011100000011010;
   assign mem[510] = 32'b11111110100101001011010000111100;
   assign mem[511] = 32'b11111010110000010010011001110000;
   assign mem[512] = 32'b00000001101000001101000010100010;
   assign mem[513] = 32'b11111011100101101000111001010000;
   assign mem[514] = 32'b11111011000110010011010011100000;
   assign mem[515] = 32'b11111011101000111111000110101000;
   assign mem[516] = 32'b00001000000101100101001000110000;
   assign mem[517] = 32'b00000011110011010001101010100100;
   assign mem[518] = 32'b00000011000011010111000110011100;
   assign mem[519] = 32'b11111010101001101100111100010000;
   assign mem[520] = 32'b11111101110010010000010111101100;
   assign mem[521] = 32'b00000101001000011101110111100000;
   assign mem[522] = 32'b00000101100101011101001101111000;
   assign mem[523] = 32'b00000100000100011011010011100000;
   assign mem[524] = 32'b11110101000110100101011110100000;
   assign mem[525] = 32'b11101111011000100100111010000000;
   assign mem[526] = 32'b00000110010101111111101101101000;
   assign mem[527] = 32'b00000011111110111000011110001000;
   assign mem[528] = 32'b11110110001100010111111111000000;
   assign mem[529] = 32'b11110010001011110010110011010000;
   assign mem[530] = 32'b11111100100101011100011111010100;
   assign mem[531] = 32'b11111000011010100100010110100000;
   assign mem[532] = 32'b00000011100100000000101100011100;
   assign mem[533] = 32'b00000000111001110111100111010011;
   assign mem[534] = 32'b11111011110000101011101011101000;
   assign mem[535] = 32'b11110111100001110001100000000000;
   assign mem[536] = 32'b00000000101100111010001110000001;
   assign mem[537] = 32'b00000010000111001111001100000000;
   assign mem[538] = 32'b00000000001111111001100000011001;
   assign mem[539] = 32'b00000010011100010000110110111100;
   assign mem[540] = 32'b11111111001011001101010110110000;
   assign mem[541] = 32'b00000001010010000100110111100110;
   assign mem[542] = 32'b00000100110010111011101010011000;
   assign mem[543] = 32'b00000110001111101101100110110000;
   assign mem[544] = 32'b11110111000010000101011001010000;
   assign mem[545] = 32'b11101000110011101001110100100000;
   assign mem[546] = 32'b11111111110001110110111011100111;
   assign mem[547] = 32'b11111101110110010110011010111000;
   assign mem[548] = 32'b11110101010101010011111011010000;
   assign mem[549] = 32'b11110110000100000010000111100000;
   assign mem[550] = 32'b11111111100111110000100111011000;
   assign mem[551] = 32'b11111000101010011010110101110000;
   assign mem[552] = 32'b11111101101101000110010100000000;
   assign mem[553] = 32'b11111011100110111000110000101000;
   assign mem[554] = 32'b11111110111110010110101101010100;
   assign mem[555] = 32'b00000000101001000111100110010100;
   assign mem[556] = 32'b00000000011011100000110001101110;
   assign mem[557] = 32'b00000100000100001010111110000000;
   assign mem[558] = 32'b00001001100000000001101101000000;
   assign mem[559] = 32'b11111110110110111000010001111000;
   assign mem[560] = 32'b11111100010000000101111000011000;
   assign mem[561] = 32'b11111110001111010000100001001000;
   assign mem[562] = 32'b11111110010100111000000101100100;
   assign mem[563] = 32'b00000101001001010100111011110000;
   assign mem[564] = 32'b00000000000101000111000000001011;
   assign mem[565] = 32'b11111111000010110001010111110110;
   assign mem[566] = 32'b00000100010111010111000011010000;
   assign mem[567] = 32'b11111101011001101100101010101000;
   assign mem[568] = 32'b00000001100000101011010011001100;
   assign mem[569] = 32'b11111001011001101010100000011000;
   assign mem[570] = 32'b11111001110001110111100001001000;
   assign mem[571] = 32'b00001000000010101100111110110000;
   assign mem[572] = 32'b11111100110011011101011100111000;
   assign mem[573] = 32'b11111110011110100000111111010110;
   assign mem[574] = 32'b00000111011010101011110011001000;
   assign mem[575] = 32'b11111001110110111000001111010000;
   assign mem[576] = 32'b00000011011010100011000010111000;
   assign mem[577] = 32'b00000110011111101111110000110000;
   assign mem[578] = 32'b00000001101010111011101001110110;
   assign mem[579] = 32'b11101011010100100110100111100000;
   assign mem[580] = 32'b00000010011111001100111101011100;
   assign mem[581] = 32'b00000001111111101011100010101110;
   assign mem[582] = 32'b00000000101010011111110110110011;
   assign mem[583] = 32'b11111111110101100000011010011000;
   assign mem[584] = 32'b11111100011010111100011001111000;
   assign mem[585] = 32'b00000000001010001111111010000011;
   assign mem[586] = 32'b11110101110101101001010101010000;
   assign mem[587] = 32'b11111111100100000000010111100101;
   assign mem[588] = 32'b00000001111011101010010001011010;
   assign mem[589] = 32'b00000001101011001010111010000000;
   assign mem[590] = 32'b11111101111000000000111111000000;
   assign mem[591] = 32'b00000010101001011110110011001000;
   assign mem[592] = 32'b11111010101100111111011010110000;
   assign mem[593] = 32'b00000000011110000001000001011110;
   assign mem[594] = 32'b11111101001000100100010110100000;
   assign mem[595] = 32'b11111011000011100011101111011000;
   assign mem[596] = 32'b00000100111110000111100110000000;
   assign mem[597] = 32'b00000111100110011110000111111000;
   assign mem[598] = 32'b00000000101110010001100110001110;
   assign mem[599] = 32'b11111101110011110111110000110100;
   assign mem[600] = 32'b00000101011000000111010000100000;
   assign mem[601] = 32'b11111100000000110001001111101000;
   assign mem[602] = 32'b11111110000110001111011110000100;
   assign mem[603] = 32'b11111100111110010010100111110100;
   assign mem[604] = 32'b00000000111110010000011001100111;
   assign mem[605] = 32'b11111010101110001000111111111000;
   assign mem[606] = 32'b11111100001110110100110100110000;
   assign mem[607] = 32'b11111111110110010100110101111000;
   assign mem[608] = 32'b00000000100110001101111000111111;
   assign mem[609] = 32'b11111011000010011010100010000000;
   assign mem[610] = 32'b11111011111110000111101011011000;
   assign mem[611] = 32'b11111000110010101011111100001000;
   assign mem[612] = 32'b11111101110101011100100000111000;
   assign mem[613] = 32'b00000110100011110110000110111000;
   assign mem[614] = 32'b00000011100100100101100000010100;
   assign mem[615] = 32'b11111010010001110100101010111000;
   assign mem[616] = 32'b00000111001001100000010100011000;
   assign mem[617] = 32'b11111011001111110101001101101000;
   assign mem[618] = 32'b00000001001100101110110011111000;
   assign mem[619] = 32'b11111010110011011110001101011000;
   assign mem[620] = 32'b00000001000111111110100011010110;
   assign mem[621] = 32'b11111110000101110011001101010110;
   assign mem[622] = 32'b11111001011000010010001010110000;
   assign mem[623] = 32'b00000001011011101001111000110010;
   assign mem[624] = 32'b11111110110001111101111000110000;
   assign mem[625] = 32'b00000001101001011100111110101110;
   assign mem[626] = 32'b00000111101100001000101000110000;
   assign mem[627] = 32'b00000001110110101111101101101010;
   assign mem[628] = 32'b00000010110000001111010001001100;
   assign mem[629] = 32'b00000001110001011101011110100010;
   assign mem[630] = 32'b00000001101010000110100111111100;
   assign mem[631] = 32'b11111011110100011100100101101000;
   assign mem[632] = 32'b00000000111101110011100110011010;
   assign mem[633] = 32'b11111001111101110101111000010000;
   assign mem[634] = 32'b11111110111100101000111100000100;
   assign mem[635] = 32'b11111011110101101111110111001000;
   assign mem[636] = 32'b00000011000011111000100011111100;
   assign mem[637] = 32'b11110111111100111111111100100000;
   assign mem[638] = 32'b11111111100110010111000100000111;
   assign mem[639] = 32'b11111110100010011010101000011010;
   assign mem[640] = 32'b11111011011110100111101110111000;
   assign mem[641] = 32'b11111100011011011011010001010000;
   assign mem[642] = 32'b00000000001010001100010000000101;
   assign mem[643] = 32'b00000011100110011111000011001000;
   assign mem[644] = 32'b11111010010000001001011100011000;
   assign mem[645] = 32'b00001010000111010010000110100000;
   assign mem[646] = 32'b11101111101100111111000000000000;
   assign mem[647] = 32'b00000110001011100011001111110000;
   assign mem[648] = 32'b11111101010000110100101100001100;
   assign mem[649] = 32'b11111101100101010110111111010000;
   assign mem[650] = 32'b11111001110000011010011010100000;
   assign mem[651] = 32'b00000100111111111010000111011000;
   assign mem[652] = 32'b11111101000001001101101001101100;
   assign mem[653] = 32'b11111110101111111000011010001000;
   assign mem[654] = 32'b00001001011011011101010100000000;
   assign mem[655] = 32'b11110001100001001011101001000000;
   assign mem[656] = 32'b00000010000100000110101101111000;
   assign mem[657] = 32'b00001000001111010101100110100000;
   assign mem[658] = 32'b11111100101001010100100011001000;
   assign mem[659] = 32'b11101100100111010010001111100000;
   assign mem[660] = 32'b11111111110110000000100010010001;
   assign mem[661] = 32'b00001010001010010010110111100000;
   assign mem[662] = 32'b00001000110100011111010011000000;
   assign mem[663] = 32'b00000001101100010000001101100010;
   assign mem[664] = 32'b11111111110000010101111010001010;
   assign mem[665] = 32'b11111010100011011000001110001000;
   assign mem[666] = 32'b11110101110001111100010101100000;
   assign mem[667] = 32'b00000001111111100101001110100000;
   assign mem[668] = 32'b11111011110000001111111000001000;
   assign mem[669] = 32'b11110101101110001101010010110000;
   assign mem[670] = 32'b11110101100100111010111110110000;
   assign mem[671] = 32'b11111101010011001110011100001000;
   assign mem[672] = 32'b00000111111010010011100110001000;
   assign mem[673] = 32'b00000101011110001100100100101000;
   assign mem[674] = 32'b11111010010111100011001110001000;
   assign mem[675] = 32'b11100111011011010010010001000000;
   assign mem[676] = 32'b11110100111110110100001111100000;
   assign mem[677] = 32'b11111100100111000110001000101100;
   assign mem[678] = 32'b11111100101110110000001111110000;
   assign mem[679] = 32'b11111101110011101111001001110000;
   assign mem[680] = 32'b00000000010111011100011000100100;
   assign mem[681] = 32'b11111001011111000101110110010000;
   assign mem[682] = 32'b00001101010110011100010000110000;
   assign mem[683] = 32'b00000101100001010010010101111000;
   assign mem[684] = 32'b11111101111010110001010110110100;
   assign mem[685] = 32'b11110100111011001000100100110000;
   assign mem[686] = 32'b11111100000000011000100111111000;
   assign mem[687] = 32'b11110111011000111110100100010000;
   assign mem[688] = 32'b00000001101010100010010111111110;
   assign mem[689] = 32'b00000100100000000100100110001000;
   assign mem[690] = 32'b11111100101011000110101010011100;
   assign mem[691] = 32'b11111011011110000101010101010000;
   assign mem[692] = 32'b11111111101100101011011000110011;
   assign mem[693] = 32'b00001000100100100100111011010000;
   assign mem[694] = 32'b11110101010010100000100101000000;
   assign mem[695] = 32'b11111100101101011011101000101000;
   assign mem[696] = 32'b00001001001110010100100010000000;
   assign mem[697] = 32'b11111101000100101010001010100100;
   assign mem[698] = 32'b11111110011001011000011010010010;
   assign mem[699] = 32'b00000000000011111000011111000100;
   assign mem[700] = 32'b00000000001111111100110011100000;
   assign mem[701] = 32'b00000110110100110010100000110000;
   assign mem[702] = 32'b11111101100111111001101110110100;
   assign mem[703] = 32'b11110011001001000101110110100000;
   assign mem[704] = 32'b11111111100010101010111111101111;
   assign mem[705] = 32'b00000111011010101101100111001000;
   assign mem[706] = 32'b00001101011101110011110010010000;
   assign mem[707] = 32'b00000001001100011110010010111100;
   assign mem[708] = 32'b11111010101110000101000101100000;
   assign mem[709] = 32'b00000000010010101100000110010010;
   assign mem[710] = 32'b11110110110111010110001001100000;
   assign mem[711] = 32'b11111000100101000100001001100000;
   assign mem[712] = 32'b00000111010000001010001011000000;
   assign mem[713] = 32'b11111110011111100000101110000000;
   assign mem[714] = 32'b00000010100111011110011001001100;
   assign mem[715] = 32'b11111101011100111010110000001000;
   assign mem[716] = 32'b00001011101010110111100011110000;
   assign mem[717] = 32'b11110011110011101010101111100000;
   assign mem[718] = 32'b00000101011100111001001000010000;
   assign mem[719] = 32'b11111001011010010001111000001000;
   assign mem[720] = 32'b11111101111100011011000100001100;
   assign mem[721] = 32'b11111100110110000101000010110000;
   assign mem[722] = 32'b11111111110110010111011100100000;
   assign mem[723] = 32'b00000010001110101000111001101000;
   assign mem[724] = 32'b00000001101000011011111100001110;
   assign mem[725] = 32'b11111111101011010100111110101001;
   assign mem[726] = 32'b11110110101010011000110011110000;
   assign mem[727] = 32'b00000001110001101111011001101110;
   assign mem[728] = 32'b11111101100111001101101110111100;
   assign mem[729] = 32'b00000001101100110011011111111000;
   assign mem[730] = 32'b11111101111111010111100000011100;
   assign mem[731] = 32'b00000101000110001110011000111000;
   assign mem[732] = 32'b11111101100100001111110000110100;
   assign mem[733] = 32'b11111001101111010110001100001000;
   assign mem[734] = 32'b00000110000001001010110000001000;
   assign mem[735] = 32'b00000010011110111011100100110000;
   assign mem[736] = 32'b00000110101000010010010111100000;
   assign mem[737] = 32'b00000111100111011110000010001000;
   assign mem[738] = 32'b00000011110111110000010011100000;
   assign mem[739] = 32'b11111111101110000111111100100101;
   assign mem[740] = 32'b11111010000101100110100000100000;
   assign mem[741] = 32'b11110101010010000011010110000000;
   assign mem[742] = 32'b00000011011101011100111111101000;
   assign mem[743] = 32'b00000110010000000100000011011000;
   assign mem[744] = 32'b11110110011010101110011000000000;
   assign mem[745] = 32'b11111110011100000101111101001000;
   assign mem[746] = 32'b11110110101011101110000001110000;
   assign mem[747] = 32'b00000001011001011111101101110100;
   assign mem[748] = 32'b00000101001101101011011110010000;
   assign mem[749] = 32'b00001000100001110011101000000000;
   assign mem[750] = 32'b11110101111100010010001100110000;
   assign mem[751] = 32'b00001001111001101001100101110000;
   assign mem[752] = 32'b00000001110010101110010100100100;
   assign mem[753] = 32'b00000110011100101101010110010000;
   assign mem[754] = 32'b11111111100101010001011110111111;
   assign mem[755] = 32'b00000001111101001011101000101000;
   assign mem[756] = 32'b11110100011000110101001101010000;
   assign mem[757] = 32'b00001011010000010011000000100000;
   assign mem[758] = 32'b11111100100000101010001111101100;
   assign mem[759] = 32'b11100010000110000110100010000000;
   assign mem[760] = 32'b11111101100111110101101110100100;
   assign mem[761] = 32'b11110110111010111000010010000000;
   assign mem[762] = 32'b11111101111100110101100011100100;
   assign mem[763] = 32'b00000100010110101011101011101000;
   assign mem[764] = 32'b11111111000110011010011101110101;
   assign mem[765] = 32'b00000101111111101001010110111000;
   assign mem[766] = 32'b11101100110011011110100001100000;
   assign mem[767] = 32'b00000010111011000110110111110000;
   assign mem[768] = 32'b11111110010000000101101101101000;
   assign mem[769] = 32'b00000001111100100010101111110100;
   assign mem[770] = 32'b11111110111011000001010000001000;
   assign mem[771] = 32'b11111100100010011010101010110000;
   assign mem[772] = 32'b00000011001010110111010100011000;
   assign mem[773] = 32'b11111111101010110101011100011011;
   assign mem[774] = 32'b11111110010010111001001000010100;
   assign mem[775] = 32'b00000001011001111000101100101000;
   assign mem[776] = 32'b11110111010110001011101100010000;
   assign mem[777] = 32'b00000011111111111000100010110100;
   assign mem[778] = 32'b11111110001101100011000101100100;
   assign mem[779] = 32'b11111111011101001101001011101011;
   assign mem[780] = 32'b00000011010001010101001101010000;
   assign mem[781] = 32'b11111101110011011111111110001000;
   assign mem[782] = 32'b11111010111101110110000001110000;
   assign mem[783] = 32'b00000010101001110110110101101000;
   assign mem[784] = 32'b11110110000011110110101010000000;
   assign mem[785] = 32'b00000011100010100001110110000000;
   assign mem[786] = 32'b11111111010001001100100100101001;
   assign mem[787] = 32'b00000111111001000110011111110000;
   assign mem[788] = 32'b11111110010101111000110011111000;
   assign mem[789] = 32'b00000011010110001000010110010100;
   assign mem[790] = 32'b00000001000010010111011111110000;
   assign mem[791] = 32'b11111011000100110111011011100000;
   assign mem[792] = 32'b11111110001100101010110110011110;
   assign mem[793] = 32'b11111001111110011110001101011000;
   assign mem[794] = 32'b00000000111110001001011000111110;
   assign mem[795] = 32'b11111011110010110100100100010000;
   assign mem[796] = 32'b00000010010100100001111010000100;
   assign mem[797] = 32'b11111101000001110101111000000000;
   assign mem[798] = 32'b00000001100100101111111010010100;
   assign mem[799] = 32'b11111110110110101001011110011010;
   assign mem[800] = 32'b11110101011101011100011111010000;
   assign mem[801] = 32'b11110110000110000001100101110000;
   assign mem[802] = 32'b11111111111011100101001100011011;
   assign mem[803] = 32'b00000000110001001011110110011010;
   assign mem[804] = 32'b00000110111110110110001111010000;
   assign mem[805] = 32'b11111101011101001111000101001000;
   assign mem[806] = 32'b11111010010100000010000000001000;
   assign mem[807] = 32'b00001100011011110010000001100000;
   assign mem[808] = 32'b11111011000110001110110101110000;
   assign mem[809] = 32'b00000011101010011110010001100000;
   assign mem[810] = 32'b00000000000111001011101100000010;
   assign mem[811] = 32'b00000000111011101000000101111010;
   assign mem[812] = 32'b00000010111011100000010111011000;
   assign mem[813] = 32'b00000101001010000110001011101000;
   assign mem[814] = 32'b11111100110101101101100000100000;
   assign mem[815] = 32'b11111101010001011000110001011100;
   assign mem[816] = 32'b00000010101100110011101011100100;
   assign mem[817] = 32'b11111011000010110000000010100000;
   assign mem[818] = 32'b00000110010111011000101100101000;
   assign mem[819] = 32'b11111011000101101010011000110000;
   assign mem[820] = 32'b00000001110111011011100101111100;
   assign mem[821] = 32'b00000010110001111011101111000000;
   assign mem[822] = 32'b11111101010000010110000000100100;
   assign mem[823] = 32'b11111110010010111000101110110110;
   assign mem[824] = 32'b00000110001110011100011101001000;
   assign mem[825] = 32'b11110100000001001111001110100000;
   assign mem[826] = 32'b11111010100110111100011011000000;
   assign mem[827] = 32'b00001100101001001010001110100000;
   assign mem[828] = 32'b11111010011000011000010111010000;
   assign mem[829] = 32'b11110011011111000010111000010000;
   assign mem[830] = 32'b00000010100001111000110000000100;
   assign mem[831] = 32'b11111010001011010011011111011000;
   assign mem[832] = 32'b11111100101110100110101101010000;
   assign mem[833] = 32'b00000010010000101001101100101100;
   assign mem[834] = 32'b00000000001010001111111110001111;
   assign mem[835] = 32'b11111111110110011100001000110100;
   assign mem[836] = 32'b11110101000001011100001010100000;
   assign mem[837] = 32'b11111101001011001101101100000000;
   assign mem[838] = 32'b00000100100110010010011111111000;
   assign mem[839] = 32'b00000000101100100000011011111101;
   assign mem[840] = 32'b11111101110100010001111010100000;
   assign mem[841] = 32'b11111111001011000001011111110010;
   assign mem[842] = 32'b00000001101001111100101111000000;
   assign mem[843] = 32'b11110110100101000100010010110000;
   assign mem[844] = 32'b00000011011001100010111111111100;
   assign mem[845] = 32'b00000101010100110011101000111000;
   assign mem[846] = 32'b00001100111000101110110110010000;
   assign mem[847] = 32'b00000010100000101111100110000000;
   assign mem[848] = 32'b11111001100011011100111100001000;
   assign mem[849] = 32'b11111110011111001001100010101110;
   assign mem[850] = 32'b11111111011100101001111101000010;
   assign mem[851] = 32'b11111000111111000110101110011000;
   assign mem[852] = 32'b11111101101110100001010101100100;
   assign mem[853] = 32'b00000010111010001010101101011000;
   assign mem[854] = 32'b11110111100001000011000100000000;
   assign mem[855] = 32'b11111101111110111111110100000000;
   assign mem[856] = 32'b11110110111010001001011111100000;
   assign mem[857] = 32'b00000000001010101111010011110110;
   assign mem[858] = 32'b00000001110011100101010101111010;
   assign mem[859] = 32'b00001000100110011111001101100000;
   assign mem[860] = 32'b11110011110010100011101000100000;
   assign mem[861] = 32'b11110010101100111111100001110000;
   assign mem[862] = 32'b00000000110001001011001010000010;
   assign mem[863] = 32'b11111110001001100000101011001110;
   assign mem[864] = 32'b00000101111111011011111011011000;
   assign mem[865] = 32'b00000000101111101000001110000011;
   assign mem[866] = 32'b00000011111011011001010111110000;
   assign mem[867] = 32'b00000001010011110111011001001000;
   assign mem[868] = 32'b00000111011100110101100111010000;
   assign mem[869] = 32'b00000010010001101101001111110100;
   assign mem[870] = 32'b11110111110101110111100101000000;
   assign mem[871] = 32'b00000111000010100000101010010000;
   assign mem[872] = 32'b11111011110101110010101110100000;
   assign mem[873] = 32'b00000101111000111000010101000000;
   assign mem[874] = 32'b11111011100011101010110101010000;
   assign mem[875] = 32'b00000111110101110101011110110000;
   assign mem[876] = 32'b00000011001011011000101100010000;
   assign mem[877] = 32'b00000110010100101101110001001000;
   assign mem[878] = 32'b11111100100000111101100011000100;
   assign mem[879] = 32'b11101011011100000011010100000000;
   assign mem[880] = 32'b11101111101011101010101111000000;
   assign mem[881] = 32'b00001011110000100111000110010000;
   assign mem[882] = 32'b00000010110101000000001101000000;
   assign mem[883] = 32'b00000010001101001111111110100100;
   assign mem[884] = 32'b00001010110001000101011011110000;
   assign mem[885] = 32'b00001010010001101100010100010000;
   assign mem[886] = 32'b00000010001011001100000101100100;
   assign mem[887] = 32'b00000111001000101000111000101000;
   assign mem[888] = 32'b11110001111111111111101001100000;
   assign mem[889] = 32'b11101011011011010110010110000000;
   assign mem[890] = 32'b11110100100001010111000010000000;
   assign mem[891] = 32'b11111111010010101111011111100000;
   assign mem[892] = 32'b11110010100101000110000010110000;
   assign mem[893] = 32'b00000111011000101011101011010000;
   assign mem[894] = 32'b00000000111000010101010000000111;
   assign mem[895] = 32'b11101111101001001011001110100000;
   assign mem[896] = 32'b00010010111001100011101010000000;
   assign mem[897] = 32'b11111001100101011001100010100000;
   assign mem[898] = 32'b11111001001100111110011011001000;
   assign mem[899] = 32'b11100111100101010000100010000000;
   assign mem[900] = 32'b11110100111010100101011010110000;
   assign mem[901] = 32'b00000101011111101100011001010000;
   assign mem[902] = 32'b11101001011010101010010010000000;
   assign mem[903] = 32'b00001111100011010101000010100000;
   assign mem[904] = 32'b00000100010001101000000010011000;
   assign mem[905] = 32'b11110100100110001000110011110000;
   assign mem[906] = 32'b00001001011100111111100010100000;
   assign mem[907] = 32'b11111110100101111100101011010100;
   assign mem[908] = 32'b11111011110101010001000000111000;
   assign mem[909] = 32'b11100100101000001011011100100000;
   assign mem[910] = 32'b11111100001011110100011001000100;
   assign mem[911] = 32'b11111011101111000111100110100000;
   assign mem[912] = 32'b00000010011100111000010110110100;
   assign mem[913] = 32'b11111110111110001110011101111110;
   assign mem[914] = 32'b00000000110111000100010111000001;
   assign mem[915] = 32'b11111101110100010111011010111000;
   assign mem[916] = 32'b11111110001101001000010001111000;
   assign mem[917] = 32'b00000010100100010011100000010100;
   assign mem[918] = 32'b00000000111101000110001101000000;
   assign mem[919] = 32'b00000100000011001001101110110000;
   assign mem[920] = 32'b00000001001000001000011101100110;
   assign mem[921] = 32'b11111000100110001001100000011000;
   assign mem[922] = 32'b11111101100001011010101110010100;
   assign mem[923] = 32'b00000011000100111001111010000100;
   assign mem[924] = 32'b11110101101010010001111000100000;
   assign mem[925] = 32'b00000111000111110000101011110000;
   assign mem[926] = 32'b11111011001011011111001100001000;
   assign mem[927] = 32'b00000001000000110110001110011110;
   assign mem[928] = 32'b00000001001100001101000111100100;
   assign mem[929] = 32'b00000111111111011101011101110000;
   assign mem[930] = 32'b00000000001110011010000000101110;
   assign mem[931] = 32'b00000000011111000100100000110111;
   assign mem[932] = 32'b11111111110010100110011110000001;
   assign mem[933] = 32'b00000010010011010101011011101100;
   assign mem[934] = 32'b11111101101000000000010100100000;
   assign mem[935] = 32'b00000010100011011000111111011100;
   assign mem[936] = 32'b11110100111100011110100000100000;
   assign mem[937] = 32'b00000010110010011111010000010100;
   assign mem[938] = 32'b00000000001100110010100010101011;
   assign mem[939] = 32'b00000000111101000101111001101010;
   assign mem[940] = 32'b11111011000010011000011011101000;
   assign mem[941] = 32'b11111110100110001000000110100000;
   assign mem[942] = 32'b11110110111001011001111110010000;
   assign mem[943] = 32'b11111010111000000110101001001000;
   assign mem[944] = 32'b00001010110111000101000010100000;
   assign mem[945] = 32'b00000111101001011101001111011000;
   assign mem[946] = 32'b00001110101101110000101110000000;
   assign mem[947] = 32'b11111010100001010010111101001000;
   assign mem[948] = 32'b11111011111100000110010100001000;
   assign mem[949] = 32'b11100001101111101100101010100000;
   assign mem[950] = 32'b11101101111011101001010100100000;
   assign mem[951] = 32'b11111101101011010011001100111100;
   assign mem[952] = 32'b00000111110001011110010101010000;
   assign mem[953] = 32'b00000000100100001110111010101000;
   assign mem[954] = 32'b00000000000001001100111000101011;
   assign mem[955] = 32'b11110101111011011110010101010000;
   assign mem[956] = 32'b11111000110110100000011101110000;
   assign mem[957] = 32'b00001011100110111000000100100000;
   assign mem[958] = 32'b11111101111100010110100100010100;
   assign mem[959] = 32'b00000001100010000000010111010100;
   assign mem[960] = 32'b11110110111111100001110010010000;
   assign mem[961] = 32'b11101111000001011001000100100000;
   assign mem[962] = 32'b00000000100000000000010101010000;
   assign mem[963] = 32'b00000000001010111001100011100010;
   assign mem[964] = 32'b00000000101110101011001000011100;
   assign mem[965] = 32'b00000100100010111010111111001000;
   assign mem[966] = 32'b00000100101010101111100000000000;
   assign mem[967] = 32'b11111110101100001100100000111100;
   assign mem[968] = 32'b00000000001101110000111010000000;
   assign mem[969] = 32'b00001011111100010000100001110000;
   assign mem[970] = 32'b00000001000100100111111101001100;
   assign mem[971] = 32'b00000000100010100000000111010001;
   assign mem[972] = 32'b00000010101000111001110100000000;
   assign mem[973] = 32'b00000010001011110101011000100000;
   assign mem[974] = 32'b11111101110100001010110111000100;
   assign mem[975] = 32'b11111011101100111100101101010000;
   assign mem[976] = 32'b00000100011010001010100100000000;
   assign mem[977] = 32'b00000011011101111110000110010000;
   assign mem[978] = 32'b00001000100010111011011011010000;
   assign mem[979] = 32'b11111100110101001110100010011100;
   assign mem[980] = 32'b11111011111111110111110001111000;
   assign mem[981] = 32'b11110010010101110111111101010000;
   assign mem[982] = 32'b00000000001100000100010110001100;
   assign mem[983] = 32'b00000100111001111100111110011000;
   assign mem[984] = 32'b11101110001110111011010010100000;
   assign mem[985] = 32'b11111100001110101111011010011000;
   assign mem[986] = 32'b00000010110110000000011101100100;
   assign mem[987] = 32'b11111111010011011110010011100100;
   assign mem[988] = 32'b00000111001111111111010001010000;
   assign mem[989] = 32'b00000101010010110000011001001000;
   assign mem[990] = 32'b11111001001001001101101011010000;
   assign mem[991] = 32'b11111110001001100011010001110100;
   assign mem[992] = 32'b11111111100011001011010011000111;
   assign mem[993] = 32'b11111100111000001100011011100100;
   assign mem[994] = 32'b11111010111101010101010110000000;
   assign mem[995] = 32'b11111110101000001000101001111010;
   assign mem[996] = 32'b11111011110100100110110110011000;
   assign mem[997] = 32'b11111101001101001010000111110100;
   assign mem[998] = 32'b00000001001110011000110100000100;
   assign mem[999] = 32'b00000110001101011101000100001000;
   assign mem[1000] = 32'b11111111011001111010110011001001;
   assign mem[1001] = 32'b00000000100010110001110011110001;
   assign mem[1002] = 32'b00000100010111010110110001010000;
   assign mem[1003] = 32'b11111111100010110000110011000010;
   assign mem[1004] = 32'b00000001111011111100101011110010;
   assign mem[1005] = 32'b00000000000110010001110001011001;
   assign mem[1006] = 32'b11110010100101100000111110000000;
   assign mem[1007] = 32'b00000110001101111000000101001000;
   assign mem[1008] = 32'b11111010001111001001111010000000;
   assign mem[1009] = 32'b11111001101100110100101001000000;
   assign mem[1010] = 32'b11111101111011000110111110101100;
   assign mem[1011] = 32'b00001000001101110001100100110000;
   assign mem[1012] = 32'b11111100010001101010011011110100;
   assign mem[1013] = 32'b00000010011001101001010101110000;
   assign mem[1014] = 32'b00001111110100010101000100110000;
   assign mem[1015] = 32'b00000010100010000001000011011000;
   assign mem[1016] = 32'b11111010010000101100100000010000;
   assign mem[1017] = 32'b00000011011111101001011010011000;
   assign mem[1018] = 32'b11111011001100010010011100110000;
   assign mem[1019] = 32'b11110010010101000101010000110000;
   assign mem[1020] = 32'b00000010000001111110001111100100;
   assign mem[1021] = 32'b11111011000101101011100100011000;
   assign mem[1022] = 32'b00000010001110011000001110111100;
   assign mem[1023] = 32'b00000010101101110000100010000000;
   assign mem[1024] = 32'b11111100011100110011110010110100;
   assign mem[1025] = 32'b11111000111101110001110001101000;
   assign mem[1026] = 32'b00001010110101011110111100100000;
   assign mem[1027] = 32'b00000010011110001110010000111100;
   assign mem[1028] = 32'b11111001001001011101000100010000;
   assign mem[1029] = 32'b11111100010100000100111010011000;
   assign mem[1030] = 32'b00000010100000100110111111000100;
   assign mem[1031] = 32'b11110110001011011001001000010000;
   assign mem[1032] = 32'b00000011100001100001110001111100;
   assign mem[1033] = 32'b00000011101000000011011000001000;
   assign mem[1034] = 32'b11111111010001010101010101111001;
   assign mem[1035] = 32'b11111101111110000000111100100100;
   assign mem[1036] = 32'b11111001001001110010110110101000;
   assign mem[1037] = 32'b00000001000000000000100100111010;
   assign mem[1038] = 32'b00000010100011011000101110111000;
   assign mem[1039] = 32'b00000000110011111100100100101010;
   assign mem[1040] = 32'b11110101101111111100011111110000;
   assign mem[1041] = 32'b11111100000100110100110111000000;
   assign mem[1042] = 32'b00001010111100000101000100110000;
   assign mem[1043] = 32'b00000111010100001110000000101000;
   assign mem[1044] = 32'b11110100000001010111000011100000;
   assign mem[1045] = 32'b11110011000110110010001011010000;
   assign mem[1046] = 32'b11111101110001011110100100001100;
   assign mem[1047] = 32'b11110111110111010101100101110000;
   assign mem[1048] = 32'b11111101111110001111010001101000;
   assign mem[1049] = 32'b11111001111100110000010100100000;
   assign mem[1050] = 32'b11110001100111110011010110000000;
   assign mem[1051] = 32'b11101101001010100001110001100000;
   assign mem[1052] = 32'b00000110100100111001110010111000;
   assign mem[1053] = 32'b00000111000111000000110010101000;
   assign mem[1054] = 32'b11110110000001101011000100010000;
   assign mem[1055] = 32'b11110010111001111001000001000000;
   assign mem[1056] = 32'b11111110101000100010100001111100;
   assign mem[1057] = 32'b11110000101001010101011101100000;
   assign mem[1058] = 32'b11111001101000011001100011100000;
   assign mem[1059] = 32'b11111100011110111010100110000000;
   assign mem[1060] = 32'b11110001100101000111101110010000;
   assign mem[1061] = 32'b11111011101101011010111001010000;
   assign mem[1062] = 32'b00001011001000010111100010010000;
   assign mem[1063] = 32'b00000111100001001010111110011000;
   assign mem[1064] = 32'b11111100111110000101000010111100;
   assign mem[1065] = 32'b11101100111000111000100101000000;
   assign mem[1066] = 32'b11111101011001000110111011111100;
   assign mem[1067] = 32'b00001001101110000001011010000000;
   assign mem[1068] = 32'b11111100000010000001000000110100;
   assign mem[1069] = 32'b11111111000001011110110000011011;
   assign mem[1070] = 32'b11111000100101011001011111100000;
   assign mem[1071] = 32'b00000101010100101111001000110000;
   assign mem[1072] = 32'b11111000001101110100011110101000;
   assign mem[1073] = 32'b00000000100010110011101010011101;
   assign mem[1074] = 32'b00001101101000101011101110110000;
   assign mem[1075] = 32'b00000010001111000011001010001000;
   assign mem[1076] = 32'b00001001001101001001001011100000;
   assign mem[1077] = 32'b11111011100110000011100001001000;
   assign mem[1078] = 32'b11110011100001111100100000100000;
   assign mem[1079] = 32'b11101001011101100011101001100000;
   assign mem[1080] = 32'b00000010110110100111000101100000;
   assign mem[1081] = 32'b11111111011011100100100100001010;
   assign mem[1082] = 32'b00000011001101111101000110011000;
   assign mem[1083] = 32'b00000111000000010010111010110000;
   assign mem[1084] = 32'b11110101010000110100010011100000;
   assign mem[1085] = 32'b11111011101100011010111100111000;
   assign mem[1086] = 32'b00000011000100001010101110001100;
   assign mem[1087] = 32'b00000011010110111000110101000100;
   assign mem[1088] = 32'b11110111011111100101111000100000;
   assign mem[1089] = 32'b11111111111011111000100101110000;
   assign mem[1090] = 32'b11111111111100010010111101001001;
   assign mem[1091] = 32'b00000000101001010100011101011101;
   assign mem[1092] = 32'b00000010111110111101000001101100;
   assign mem[1093] = 32'b11111011011010001011101110010000;
   assign mem[1094] = 32'b00000100111101111011001111011000;
   assign mem[1095] = 32'b11111111100001100100110001100111;
   assign mem[1096] = 32'b00000000010011011111111010010001;
   assign mem[1097] = 32'b11111111011001010101000011011101;
   assign mem[1098] = 32'b11111101101000111000010010000100;
   assign mem[1099] = 32'b11111101001110001011101011001000;
   assign mem[1100] = 32'b11111010000110001011111101010000;
   assign mem[1101] = 32'b00001010110001000000110000000000;
   assign mem[1102] = 32'b11111111010010010001101110010100;
   assign mem[1103] = 32'b11110111100000010000010011100000;
   assign mem[1104] = 32'b00000110001111111111000011100000;
   assign mem[1105] = 32'b00001110010110000100000110100000;
   assign mem[1106] = 32'b00000001010011001101101010011010;
   assign mem[1107] = 32'b11111011011111001101001010111000;
   assign mem[1108] = 32'b11111101110100000101100101110100;
   assign mem[1109] = 32'b11111001000100110011101101010000;
   assign mem[1110] = 32'b11111111101111011101011001011000;
   assign mem[1111] = 32'b11111111110000110011010110001011;
   assign mem[1112] = 32'b11111110010010100100001110010000;
   assign mem[1113] = 32'b00000010010000010000011001010100;
   assign mem[1114] = 32'b00000001111101001111001000010010;
   assign mem[1115] = 32'b11111100101100100101111101100100;
   assign mem[1116] = 32'b00000000010001111100111100011001;
   assign mem[1117] = 32'b00000001011011100100110010001110;
   assign mem[1118] = 32'b00000000111100011011001001001001;
   assign mem[1119] = 32'b00000001010011110111111011011010;
   assign mem[1120] = 32'b00000110101110001001010111000000;
   assign mem[1121] = 32'b11101110001010100001111100100000;
   assign mem[1122] = 32'b00000111100011110110101011011000;
   assign mem[1123] = 32'b11111010001110100111110000010000;
   assign mem[1124] = 32'b11110110100100111101001100110000;
   assign mem[1125] = 32'b11111100011001111110011110110100;
   assign mem[1126] = 32'b00001000100011011011000010110000;
   assign mem[1127] = 32'b11111100101010011001000010101000;
   assign mem[1128] = 32'b11111111000010001100111110001001;
   assign mem[1129] = 32'b00000000000101011010010101100000;
   assign mem[1130] = 32'b00000001001000010111101010000110;
   assign mem[1131] = 32'b11111101100011001100001110111100;
   assign mem[1132] = 32'b00000100001010010000110111011000;
   assign mem[1133] = 32'b11111011111110101000000101001000;
   assign mem[1134] = 32'b00000000111110010110001110010010;
   assign mem[1135] = 32'b11111111110111111011101110011000;
   assign mem[1136] = 32'b11111111011100101010001100010101;
   assign mem[1137] = 32'b11111101110000110110010011010000;
   assign mem[1138] = 32'b00000101000000000110000001000000;
   assign mem[1139] = 32'b11111110001100011010001110010010;
   assign mem[1140] = 32'b11111101111111110011011110000000;
   assign mem[1141] = 32'b11111111000101010010011111110111;
   assign mem[1142] = 32'b00000000010110111000100001110100;
   assign mem[1143] = 32'b00000010010111000010100000101000;
   assign mem[1144] = 32'b11110111001110000001010101010000;
   assign mem[1145] = 32'b11111000011001011101100011110000;
   assign mem[1146] = 32'b00000101110001111011001111011000;
   assign mem[1147] = 32'b11111011010001111000011101010000;
   assign mem[1148] = 32'b00001010100111011111000000110000;
   assign mem[1149] = 32'b00001011010110111001110001010000;
   assign mem[1150] = 32'b11110111001010001111110001100000;
   assign mem[1151] = 32'b00000011010001001000010000111000;
   assign mem[1152] = 32'b11111101110010000011000010100100;
   assign mem[1153] = 32'b00000010010111011000111111011000;
   assign mem[1154] = 32'b00000110000111100101011011000000;
   assign mem[1155] = 32'b11111110111100010110011110000010;
   assign mem[1156] = 32'b11111010110011001111111010000000;
   assign mem[1157] = 32'b00000000001000110011100111101111;
   assign mem[1158] = 32'b00000110110010010101001101000000;
   assign mem[1159] = 32'b11111110001100000100011101110000;
   assign mem[1160] = 32'b11110010111111110000100101100000;
   assign mem[1161] = 32'b11111111000110001101100001100100;
   assign mem[1162] = 32'b00000000111100110000110001101110;
   assign mem[1163] = 32'b00000011111001010010000100111000;
   assign mem[1164] = 32'b11111010011111100011001011000000;
   assign mem[1165] = 32'b11111110001101110110111010000010;
   assign mem[1166] = 32'b11111101011101111001100011111100;
   assign mem[1167] = 32'b00000111100000100111101000101000;
   assign mem[1168] = 32'b00000011110010010000010010110100;
   assign mem[1169] = 32'b00000000010111010111111000110101;
   assign mem[1170] = 32'b00000000111011100111110000000100;
   assign mem[1171] = 32'b11110101101011111101100100000000;
   assign mem[1172] = 32'b00000011011000010111001001000100;
   assign mem[1173] = 32'b00000000111100111110111011100000;
   assign mem[1174] = 32'b11110100000001111111010111110000;
   assign mem[1175] = 32'b00000100000110010000100011000000;
   assign mem[1176] = 32'b00000010011011011100010111001100;
   assign mem[1177] = 32'b00000100100011000010100111110000;
   assign mem[1178] = 32'b00000000001010010000001101101001;
   assign mem[1179] = 32'b00000001100100001110010001100110;
   assign mem[1180] = 32'b11110101010001111111100111000000;
   assign mem[1181] = 32'b11110100111010001110101010100000;
   assign mem[1182] = 32'b00001000011110010110111100010000;
   assign mem[1183] = 32'b00000011011001111000100010000100;
   assign mem[1184] = 32'b11110101000111010111001100100000;
   assign mem[1185] = 32'b11111110111110010111111100011100;
   assign mem[1186] = 32'b00000011011100001100111101100100;
   assign mem[1187] = 32'b00000010001110011101111100011100;
   assign mem[1188] = 32'b11111110101111011011010001011100;
   assign mem[1189] = 32'b00000101111010001100111010001000;
   assign mem[1190] = 32'b11111011011011110110001100110000;
   assign mem[1191] = 32'b00000010111101111111101010011100;
   assign mem[1192] = 32'b11111011000010101011101101111000;
   assign mem[1193] = 32'b11111101011001001001111001101000;
   assign mem[1194] = 32'b00000011010101101101111101011000;
   assign mem[1195] = 32'b00000111011000010111100110110000;
   assign mem[1196] = 32'b00001010101000101010010110100000;
   assign mem[1197] = 32'b11111101010001101111100011100000;
   assign mem[1198] = 32'b11111100010101010111100100110000;
   assign mem[1199] = 32'b11110101011000101101111000010000;
   assign mem[1200] = 32'b11110111111111000010101100010000;
   assign mem[1201] = 32'b11111111000100100110011100000100;
   assign mem[1202] = 32'b11111110001110010001111111101000;
   assign mem[1203] = 32'b11111111000111011010110011100000;
   assign mem[1204] = 32'b00000010100010110111110000011000;
   assign mem[1205] = 32'b11111001011110100110111010110000;
   assign mem[1206] = 32'b11111111100101011101110111010111;
   assign mem[1207] = 32'b11111111111100010110110000001011;
   assign mem[1208] = 32'b00001000011001010111111101110000;
   assign mem[1209] = 32'b11110100111100001101101010110000;
   assign mem[1210] = 32'b11111001111111110111011000001000;
   assign mem[1211] = 32'b00000010100011110010000000010000;
   assign mem[1212] = 32'b00000101111011001000111000101000;
   assign mem[1213] = 32'b00001001011100011011100111100000;
   assign mem[1214] = 32'b11111011110111100101011001111000;
   assign mem[1215] = 32'b11110110111010000110000110000000;
   assign mem[1216] = 32'b11111100011000101101111110100100;
   assign mem[1217] = 32'b00000101000001000110111001100000;
   assign mem[1218] = 32'b11111011000101011000001100101000;
   assign mem[1219] = 32'b11101001001101001001110101000000;
   assign mem[1220] = 32'b11111011110111110101110110010000;
   assign mem[1221] = 32'b11111100110100001001100011100100;
   assign mem[1222] = 32'b00000000111010000111110101110110;
   assign mem[1223] = 32'b00000001011000000011101111111010;
   assign mem[1224] = 32'b11111111111001000011111110010010;
   assign mem[1225] = 32'b11111011100001011010011000110000;
   assign mem[1226] = 32'b11111100001011000110011111111000;
   assign mem[1227] = 32'b00000010111100001001011110111000;
   assign mem[1228] = 32'b00000011010111011111111001111100;
   assign mem[1229] = 32'b00000001000010011100100110000100;
   assign mem[1230] = 32'b11111011010101111000000111000000;
   assign mem[1231] = 32'b00000001010110101101000101101100;
   assign mem[1232] = 32'b11111111001011110011101100011001;
   assign mem[1233] = 32'b11111110111001001000101000101110;
   assign mem[1234] = 32'b11111110100100110011001000011100;
   assign mem[1235] = 32'b00000011100110001110101010110100;
   assign mem[1236] = 32'b00000000101111101100011000110101;
   assign mem[1237] = 32'b00000011010110101000001111111000;
   assign mem[1238] = 32'b00000000010010011101100100001100;
   assign mem[1239] = 32'b11111111101111100010001011010010;
   assign mem[1240] = 32'b00000000010110010100000001101000;
   assign mem[1241] = 32'b11111101011101010111111011101000;
   assign mem[1242] = 32'b11111111011000010100111011100000;
   assign mem[1243] = 32'b00000000011001100110000110111010;
   assign mem[1244] = 32'b00000000100000000111110001011101;
   assign mem[1245] = 32'b11111111100111101101100111101011;
   assign mem[1246] = 32'b11110111111001000000011001110000;
   assign mem[1247] = 32'b11111110110000101101011010100010;
   assign mem[1248] = 32'b00000000100000101010000101100010;
   assign mem[1249] = 32'b11111101101000101100001000011100;
   assign mem[1250] = 32'b11111101011101011100111101001000;
   assign mem[1251] = 32'b11111011111000100001001001111000;
   assign mem[1252] = 32'b00000001101110100011011111010110;
   assign mem[1253] = 32'b11111111001110010000000000110000;
   assign mem[1254] = 32'b11111110101101010100101110101000;
   assign mem[1255] = 32'b11111100110110110011111101011000;
   assign mem[1256] = 32'b00000001001101000100110100101100;
   assign mem[1257] = 32'b11111100000010011010000000100100;
   assign mem[1258] = 32'b00000111011110001011111001010000;
   assign mem[1259] = 32'b11111111000111010100100001001011;
   assign mem[1260] = 32'b11111111000000101101100101111001;
   assign mem[1261] = 32'b00000100110000000101100011110000;
   assign mem[1262] = 32'b00000001001111110100011100011100;
   assign mem[1263] = 32'b11111011100000000010011101011000;
   assign mem[1264] = 32'b00000011100011110000010011110000;
   assign mem[1265] = 32'b00000000101010011001111010111011;
   assign mem[1266] = 32'b00000000001011000110100010111001;
   assign mem[1267] = 32'b00000000001000111110011100000010;
   assign mem[1268] = 32'b00000100011001100101101101111000;
   assign mem[1269] = 32'b11111101011010010000011010000000;
   assign mem[1270] = 32'b11111111100010001001110100011100;
   assign mem[1271] = 32'b00000110010101101111111000110000;
   assign mem[1272] = 32'b11111100000101111000000110110000;
   assign mem[1273] = 32'b11110110011011000010111100010000;
   assign mem[1274] = 32'b00000010101010100011100100001100;
   assign mem[1275] = 32'b00000011110000000111011111111100;
   assign mem[1276] = 32'b00000110001000001101111010011000;
   assign mem[1277] = 32'b00000011010011011100000101010000;
   assign mem[1278] = 32'b11111100110001101110100100101100;
   assign mem[1279] = 32'b11111011100111000011000011010000;
   assign mem[1280] = 32'b11111001011101100101010110101000;
   assign mem[1281] = 32'b11101111110001010000011001000000;
   assign mem[1282] = 32'b00000010000000100010110001000100;
   assign mem[1283] = 32'b00000101010100000010011111010000;
   assign mem[1284] = 32'b11111011001011110010111100101000;
   assign mem[1285] = 32'b00000011010001111101100100101000;
   assign mem[1286] = 32'b11110011000101100101100101000000;
   assign mem[1287] = 32'b00000011101011000110011101110000;
   assign mem[1288] = 32'b11111110011010001100101000011110;
   assign mem[1289] = 32'b00000000101100010110100100001111;
   assign mem[1290] = 32'b11111010110001000100010010100000;
   assign mem[1291] = 32'b00000010011110101110010100100100;
   assign mem[1292] = 32'b00000011110010011001100001011000;
   assign mem[1293] = 32'b00000010111010100100111011101100;
   assign mem[1294] = 32'b00001001111011110001011100100000;
   assign mem[1295] = 32'b11110010101011110110110010110000;
   assign mem[1296] = 32'b00000000010110000100010100001100;
   assign mem[1297] = 32'b00000101101000100011011000111000;
   assign mem[1298] = 32'b11110111110100110101000111110000;
   assign mem[1299] = 32'b11110111011101101010011000110000;
   assign mem[1300] = 32'b00000100111000001100010100111000;
   assign mem[1301] = 32'b11110111110011011110011011110000;
   assign mem[1302] = 32'b00000110111000011101100000011000;
   assign mem[1303] = 32'b00000000010101000001001100101011;
   assign mem[1304] = 32'b11110101000111100001010100110000;
   assign mem[1305] = 32'b11111000001110110011010011100000;
   assign mem[1306] = 32'b11111111001010011000001110001110;
   assign mem[1307] = 32'b11111111011110110101101100101100;
   assign mem[1308] = 32'b00000011110110101101011111011100;
   assign mem[1309] = 32'b00000101101110001011110001101000;
   assign mem[1310] = 32'b11111000001001100101010001101000;
   assign mem[1311] = 32'b11111011110111000010001011111000;
   assign mem[1312] = 32'b00000010000011000100010110100100;
   assign mem[1313] = 32'b00001011111101100111000010010000;
   assign mem[1314] = 32'b11110111111110100000011101010000;
   assign mem[1315] = 32'b11110011000101111011111100100000;
   assign mem[1316] = 32'b11111010110010010110101100110000;
   assign mem[1317] = 32'b00000010011000011101101100001000;
   assign mem[1318] = 32'b11111101011101101000010011010100;
   assign mem[1319] = 32'b00000101110110101101101100000000;
   assign mem[1320] = 32'b00000101001011100100100010111000;
   assign mem[1321] = 32'b11111000001001101110000000111000;
   assign mem[1322] = 32'b00000011101010000110111110001100;
   assign mem[1323] = 32'b00000010000000000101001001110000;
   assign mem[1324] = 32'b11101110001010010010010101000000;
   assign mem[1325] = 32'b11111001000100000011010001001000;
   assign mem[1326] = 32'b00000001100001011101011110010010;
   assign mem[1327] = 32'b11110011111111001100110111010000;
   assign mem[1328] = 32'b11111100010011101110011101100000;
   assign mem[1329] = 32'b00000100100111100000011001001000;
   assign mem[1330] = 32'b00000111010011000110010111000000;
   assign mem[1331] = 32'b00000111111000000010100101110000;
   assign mem[1332] = 32'b11111011111101100001110111010000;
   assign mem[1333] = 32'b11111100100101111100000010111100;
   assign mem[1334] = 32'b11111001010001111010111000110000;
   assign mem[1335] = 32'b11111110001001001111010011000110;
   assign mem[1336] = 32'b11111110110100111111000101111110;
   assign mem[1337] = 32'b00000001110010010110001110111000;
   assign mem[1338] = 32'b00000011111011010000101000101100;
   assign mem[1339] = 32'b00000011111001010111101111010100;
   assign mem[1340] = 32'b11101111100101101100010011100000;
   assign mem[1341] = 32'b00001101011001010001110110000000;
   assign mem[1342] = 32'b11110110001101001010001010110000;
   assign mem[1343] = 32'b11110000010000101100100111010000;
   assign mem[1344] = 32'b00001010011111001100001000000000;
   assign mem[1345] = 32'b11111101100000110101011101010000;
   assign mem[1346] = 32'b00011010000110100011110000000000;
   assign mem[1347] = 32'b11101101100010111001010101100000;
   assign mem[1348] = 32'b11111100011110111110001100001000;
   assign mem[1349] = 32'b11101001100100011011110000100000;
   assign mem[1350] = 32'b11111111001000101010110000111000;
   assign mem[1351] = 32'b00001010010010010100110110110000;
   assign mem[1352] = 32'b11111011101010101011010101101000;
   assign mem[1353] = 32'b11111010100100101011011101100000;
   assign mem[1354] = 32'b00000000000101011011110100001011;
   assign mem[1355] = 32'b00000100100111111000011011011000;
   assign mem[1356] = 32'b00000011000000011011110000011000;
   assign mem[1357] = 32'b11101000001110001111011101000000;
   assign mem[1358] = 32'b00000111010011111110010000000000;
   assign mem[1359] = 32'b11111010011110111100010111010000;
   assign mem[1360] = 32'b00000100011011011110000001011000;
   assign mem[1361] = 32'b00000000111001001011100101111000;
   assign mem[1362] = 32'b11111111101100110000111001010010;
   assign mem[1363] = 32'b00000001010010010101011101001100;
   assign mem[1364] = 32'b00000001011010010101100001001000;
   assign mem[1365] = 32'b11111101110111111101100011000100;
   assign mem[1366] = 32'b11111000011100100111101000011000;
   assign mem[1367] = 32'b00000011101100010110010000001100;
   assign mem[1368] = 32'b00000000111000100000010010011100;
   assign mem[1369] = 32'b00000010111110100001011101001100;
   assign mem[1370] = 32'b11111111001101101001011101000010;
   assign mem[1371] = 32'b00000011011010000111001001010100;
   assign mem[1372] = 32'b11111011010101011100011100110000;
   assign mem[1373] = 32'b11111001110010110110110000010000;
   assign mem[1374] = 32'b00001000110000001100100000010000;
   assign mem[1375] = 32'b00000010101100010110011011000000;
   assign mem[1376] = 32'b00000110000100100111000001011000;
   assign mem[1377] = 32'b11110010000011011011011101100000;
   assign mem[1378] = 32'b11111010000110101101001111111000;
   assign mem[1379] = 32'b11111000010011111100010110110000;
   assign mem[1380] = 32'b11111001011111110010110101111000;
   assign mem[1381] = 32'b11110110100010110011001111010000;
   assign mem[1382] = 32'b11111111010100111110010000101100;
   assign mem[1383] = 32'b00000001011100111111101010001100;
   assign mem[1384] = 32'b11110111101000011101111100010000;
   assign mem[1385] = 32'b11111110111011010001011110010110;
   assign mem[1386] = 32'b11111101010011011100010100111100;
   assign mem[1387] = 32'b00000000101111001110101101001000;
   assign mem[1388] = 32'b00000010011111101100100010010000;
   assign mem[1389] = 32'b00000011010110111101111111110000;
   assign mem[1390] = 32'b11111001101111101100000011011000;
   assign mem[1391] = 32'b00000110110001001011011001001000;
   assign mem[1392] = 32'b00000011101010001001000110011000;
   assign mem[1393] = 32'b00000100010001100010101110010000;
   assign mem[1394] = 32'b00000001110110001000100011110000;
   assign mem[1395] = 32'b11110011101101010101000101010000;
   assign mem[1396] = 32'b11111111000110101010001001110000;
   assign mem[1397] = 32'b11111110101101000011000111011110;
   assign mem[1398] = 32'b00000100000100011000000110011000;
   assign mem[1399] = 32'b11110011100100010011111111010000;
   assign mem[1400] = 32'b11111110000100110110011101110100;
   assign mem[1401] = 32'b11111011111010011000101000111000;
   assign mem[1402] = 32'b00000000111000111011011110111011;
   assign mem[1403] = 32'b00000010011011011001000100001100;
   assign mem[1404] = 32'b11110010110000101001100011000000;
   assign mem[1405] = 32'b00000000111110011011001010011100;
   assign mem[1406] = 32'b11111000000101001100011110111000;
   assign mem[1407] = 32'b00000001001010010000011100001100;
   assign mem[1408] = 32'b00000000101110010110011010100000;
   assign mem[1409] = 32'b00000010010110010011001010011000;
   assign mem[1410] = 32'b11111111000010011111010110110010;
   assign mem[1411] = 32'b11111010110100110110010100011000;
   assign mem[1412] = 32'b11111111100011100101100101011011;
   assign mem[1413] = 32'b00000000001011110010100000000011;
   assign mem[1414] = 32'b11111001011100110100110100010000;
   assign mem[1415] = 32'b11111100110110100111000000011000;
   assign mem[1416] = 32'b11110101101101101110111000000000;
   assign mem[1417] = 32'b00000011110000010100000100001000;
   assign mem[1418] = 32'b00000000000111000000010101011100;
   assign mem[1419] = 32'b00000011101110011101011111010100;
   assign mem[1420] = 32'b00000001001101011111010101010110;
   assign mem[1421] = 32'b11110111011011001010001101110000;
   assign mem[1422] = 32'b00000000100010000100101111010111;
   assign mem[1423] = 32'b00000100100000011011111110010000;
   assign mem[1424] = 32'b11110010111111100001001100010000;
   assign mem[1425] = 32'b00000100100101100011011100011000;
   assign mem[1426] = 32'b11111001011100110001000001111000;
   assign mem[1427] = 32'b00000110000001110110110011000000;
   assign mem[1428] = 32'b11111100100110101110001101000000;
   assign mem[1429] = 32'b11111010011101000101111001000000;
   assign mem[1430] = 32'b00000001000000000001010100111110;
   assign mem[1431] = 32'b00000000110111010001100001111100;
   assign mem[1432] = 32'b11111110000011001111101011001110;
   assign mem[1433] = 32'b11111011010101110100010100100000;
   assign mem[1434] = 32'b00000000011100100011111010010101;
   assign mem[1435] = 32'b00000011110011101110000110111100;
   assign mem[1436] = 32'b00000100010101010110011010011000;
   assign mem[1437] = 32'b11110101111100101000000100110000;
   assign mem[1438] = 32'b11111111110011011000111101100011;
   assign mem[1439] = 32'b11111110110001101101000101111100;
   assign mem[1440] = 32'b11111101110011010111011110100100;
   assign mem[1441] = 32'b00000000100101110000000110001101;
   assign mem[1442] = 32'b11111110111000010111000011001000;
   assign mem[1443] = 32'b11111111001010000001101100100101;
   assign mem[1444] = 32'b11110100110000111101110000100000;
   assign mem[1445] = 32'b00000110001010011001000000100000;
   assign mem[1446] = 32'b11111001100001100010001001100000;
   assign mem[1447] = 32'b00000011010100000011110010111000;
   assign mem[1448] = 32'b11111110110001000001100010100010;
   assign mem[1449] = 32'b11111110001010101001100011111010;
   assign mem[1450] = 32'b11111001000100111011011110111000;
   assign mem[1451] = 32'b11111101100100100011011011110100;
   assign mem[1452] = 32'b00000011010000111111000000111000;
   assign mem[1453] = 32'b00000000011011000011100001001101;
   assign mem[1454] = 32'b11110110000101101111111100100000;
   assign mem[1455] = 32'b11111110000101110011110010110010;
   assign mem[1456] = 32'b11110111100010001100101010010000;
   assign mem[1457] = 32'b11111110100111000101100000000010;
   assign mem[1458] = 32'b00000010111011011000011001000000;
   assign mem[1459] = 32'b00000010111100110111100101010100;
   assign mem[1460] = 32'b11111110110010101011101100101000;
   assign mem[1461] = 32'b11111101010110100001101111001100;
   assign mem[1462] = 32'b00000100010001100010101011101000;
   assign mem[1463] = 32'b00000100010000000010000111101000;
   assign mem[1464] = 32'b00000111000001000111100001110000;
   assign mem[1465] = 32'b00000000100110011011011110010110;
   assign mem[1466] = 32'b11110101001001101010101100110000;
   assign mem[1467] = 32'b00000110001000001100111110110000;
   assign mem[1468] = 32'b11111000000111101101101000100000;
   assign mem[1469] = 32'b11111110000100111101101010011110;
   assign mem[1470] = 32'b11111101100110110010111011000000;
   assign mem[1471] = 32'b00000001100000110100001010100100;
   assign mem[1472] = 32'b00000100101100110111000110110000;
   assign mem[1473] = 32'b00000001101111100010010000011010;
   assign mem[1474] = 32'b11111010100011101100010111111000;
   assign mem[1475] = 32'b00000001001011110100111011111110;
   assign mem[1476] = 32'b11111010111110111110011001101000;
   assign mem[1477] = 32'b11111110011111001001001010101010;
   assign mem[1478] = 32'b00000010011111001011000011101000;
   assign mem[1479] = 32'b00001000111010100101011010100000;
   assign mem[1480] = 32'b11111010011011001011001011001000;
   assign mem[1481] = 32'b00000101010001101011100000010000;
   assign mem[1482] = 32'b11111010001100100101111101011000;
   assign mem[1483] = 32'b11110110100101011101111110100000;
   assign mem[1484] = 32'b00000100101101100111001100001000;
   assign mem[1485] = 32'b00001000011100111111110010100000;
   assign mem[1486] = 32'b00000100100011110110000111001000;
   assign mem[1487] = 32'b11111000111001001001000101111000;
   assign mem[1488] = 32'b00000001011100001011110011101100;
   assign mem[1489] = 32'b11110101000111101001001101100000;
   assign mem[1490] = 32'b11111011100000001100111110010000;
   assign mem[1491] = 32'b11111001111011101100111001000000;
   assign mem[1492] = 32'b11111111001001001111100110010101;
   assign mem[1493] = 32'b00000001101001111110010010010100;
   assign mem[1494] = 32'b11110111111110000111110111100000;
   assign mem[1495] = 32'b11111110100001100000111101000000;
   assign mem[1496] = 32'b11111111111000000100101100100001;
   assign mem[1497] = 32'b00000000011100000000001110000110;
   assign mem[1498] = 32'b00000001111000010100110011110010;
   assign mem[1499] = 32'b00000110101000101011000001001000;
   assign mem[1500] = 32'b00000001000011001001010110100010;
   assign mem[1501] = 32'b00000100001111111001011101001000;
   assign mem[1502] = 32'b00000001010111111111101001001010;
   assign mem[1503] = 32'b11110110000011101101110011010000;
   assign mem[1504] = 32'b00000100100000111111100011111000;
   assign mem[1505] = 32'b11111111011110001000001010000010;
   assign mem[1506] = 32'b11111110010011010001010001101100;
   assign mem[1507] = 32'b11110100110110100001000010000000;
   assign mem[1508] = 32'b11111111111100101001110111110101;
   assign mem[1509] = 32'b00000001100101100000011011001110;
   assign mem[1510] = 32'b11111111110001100101011000100001;
   assign mem[1511] = 32'b00000101010010010100001000111000;
   assign mem[1512] = 32'b00000101110111110110000010010000;
   assign mem[1513] = 32'b00000000001000101001110000101001;
   assign mem[1514] = 32'b00000100001101010001101100001000;
   assign mem[1515] = 32'b11111111100001101001001101000011;
   assign mem[1516] = 32'b11111100000101111110100101100100;
   assign mem[1517] = 32'b00000101101010001011111000000000;
   assign mem[1518] = 32'b11111000110101110101101001010000;
   assign mem[1519] = 32'b11110010010111001111110001110000;
   assign mem[1520] = 32'b11111101101101101111011001001000;
   assign mem[1521] = 32'b00001100101010111100010100000000;
   assign mem[1522] = 32'b00000010011000101100001011000000;
   assign mem[1523] = 32'b11111110110000001110001010001110;
   assign mem[1524] = 32'b00000101110111010000000110111000;
   assign mem[1525] = 32'b00000000101110001010101100011010;
   assign mem[1526] = 32'b11111110001010000011111101010010;
   assign mem[1527] = 32'b11111110111001000101101100010110;
   assign mem[1528] = 32'b11111101010100001010011110001100;
   assign mem[1529] = 32'b11110010111000000110111100010000;
   assign mem[1530] = 32'b11110110111001111111010000010000;
   assign mem[1531] = 32'b00001100101001000110111000100000;
   assign mem[1532] = 32'b00000001011101101011101011100110;
   assign mem[1533] = 32'b00001010011010100110000111010000;
   assign mem[1534] = 32'b00001001111111111100111010010000;
   assign mem[1535] = 32'b11101001000000110101101100000000;
   assign mem[1536] = 32'b00001110110110001011001101110000;
   assign mem[1537] = 32'b11101001101111111000110110100000;
   assign mem[1538] = 32'b11111100011100000111010110100100;
   assign mem[1539] = 32'b11100101100000101110100111100000;
   assign mem[1540] = 32'b11110100111111000011110100110000;
   assign mem[1541] = 32'b00001011111000110000010100100000;
   assign mem[1542] = 32'b11111110011111001111010010111010;
   assign mem[1543] = 32'b11111111111101001000101011010100;
   assign mem[1544] = 32'b00001000100101100010001101000000;
   assign mem[1545] = 32'b11111100111010001111100101110100;
   assign mem[1546] = 32'b00001001000011110001100000010000;
   assign mem[1547] = 32'b00000110000000010101101010101000;
   assign mem[1548] = 32'b11110100001111101100010011110000;
   assign mem[1549] = 32'b11100110100110001110000100000000;
   assign mem[1550] = 32'b00000011011110100111011101000000;
   assign mem[1551] = 32'b00000100110101011110011001010000;
   assign mem[1552] = 32'b11111110101101000100001100101000;
   assign mem[1553] = 32'b11111100001110111001001111011000;
   assign mem[1554] = 32'b00000000010100100110101110011010;
   assign mem[1555] = 32'b00000000101000001111100101111100;
   assign mem[1556] = 32'b00000100001001000101110000110000;
   assign mem[1557] = 32'b11111110000010011111001000000110;
   assign mem[1558] = 32'b00000001110110001111100000001010;
   assign mem[1559] = 32'b00000000011001011101100011110011;
   assign mem[1560] = 32'b11111011011000011010100011100000;
   assign mem[1561] = 32'b11111101101001010101000111000100;
   assign mem[1562] = 32'b11111110011011100011010011110110;
   assign mem[1563] = 32'b00000001001011101111110011011000;
   assign mem[1564] = 32'b11110011000001010001101100010000;
   assign mem[1565] = 32'b00000100101011011110011011111000;
   assign mem[1566] = 32'b11110111111101101001000010010000;
   assign mem[1567] = 32'b00000101010000011111000111101000;
   assign mem[1568] = 32'b11111111100111010011001110000010;
   assign mem[1569] = 32'b00000010110110111001001011001100;
   assign mem[1570] = 32'b11111111011110010101011101010110;
   assign mem[1571] = 32'b11111101000001110011001100100000;
   assign mem[1572] = 32'b00000010110101111110010100011100;
   assign mem[1573] = 32'b00000100100101100110001001001000;
   assign mem[1574] = 32'b11111100100001000101001000111000;
   assign mem[1575] = 32'b00000001110000101001111010000110;
   assign mem[1576] = 32'b11111001111101111010111000011000;
   assign mem[1577] = 32'b00000010111010011100111101011100;
   assign mem[1578] = 32'b00000011010000010100111001101100;
   assign mem[1579] = 32'b00000011010111110000010010001100;
   assign mem[1580] = 32'b11110111010001100011011101010000;
   assign mem[1581] = 32'b00010000010000001000100101000000;
   assign mem[1582] = 32'b11110111110000110111010001000000;
   assign mem[1583] = 32'b11110111100101001101011010000000;
   assign mem[1584] = 32'b00010001001010101101010001000000;
   assign mem[1585] = 32'b00000111011101100110110100001000;
   assign mem[1586] = 32'b00001101100100110100011110110000;
   assign mem[1587] = 32'b00000111010100010100100111010000;
   assign mem[1588] = 32'b11110100010110011010110010000000;
   assign mem[1589] = 32'b11101000000010111111011110100000;
   assign mem[1590] = 32'b11111110001111110110101101110000;
   assign mem[1591] = 32'b11111101100011000000111100000100;
   assign mem[1592] = 32'b00000001101000101011010100111010;
   assign mem[1593] = 32'b00000000000101011111001001001010;
   assign mem[1594] = 32'b11101001101000000000101100000000;
   assign mem[1595] = 32'b00000010111011011110000100001100;
   assign mem[1596] = 32'b11111000000111100111011011010000;
   assign mem[1597] = 32'b00001001000000001100001011000000;
   assign mem[1598] = 32'b00000010000110000000011100110100;
   assign mem[1599] = 32'b00000000111110001000111001010001;
   assign mem[1600] = 32'b00000010011110110010101001111000;
   assign mem[1601] = 32'b00001001011110001111011111110000;
   assign mem[1602] = 32'b00000010100010110010000101010000;
   assign mem[1603] = 32'b00000001000011111101111100001000;
   assign mem[1604] = 32'b11111001111110001001010110001000;
   assign mem[1605] = 32'b00000011101110101101101000001000;
   assign mem[1606] = 32'b11111111111011100000110111011100;
   assign mem[1607] = 32'b11111001100001010110001110001000;
   assign mem[1608] = 32'b11111110101100010000101001101000;
   assign mem[1609] = 32'b11110111101111001100010111000000;
   assign mem[1610] = 32'b11111101110010001000110111010100;
   assign mem[1611] = 32'b00000011000100100101100000000100;
   assign mem[1612] = 32'b00000001000111110001110000110000;
   assign mem[1613] = 32'b11111101000111111111000000101000;
   assign mem[1614] = 32'b00001010010011101000010111000000;
   assign mem[1615] = 32'b00000000100001001101000011111000;
   assign mem[1616] = 32'b00000010101101001101101001000000;
   assign mem[1617] = 32'b11110001001101010100110011100000;
   assign mem[1618] = 32'b11111111011100000101100100010001;
   assign mem[1619] = 32'b11111011100011110001000101000000;
   assign mem[1620] = 32'b00000000011100000100000110000100;
   assign mem[1621] = 32'b11111000000101000010110111101000;
   assign mem[1622] = 32'b00000001011101110010000011010000;
   assign mem[1623] = 32'b00000011001100001011010000001000;
   assign mem[1624] = 32'b11101011111011101001001011000000;
   assign mem[1625] = 32'b00000101100111001010001011001000;
   assign mem[1626] = 32'b11111111011111110001101011001100;
   assign mem[1627] = 32'b00000010011101001001000100001100;
   assign mem[1628] = 32'b00000010110000010001110100110100;
   assign mem[1629] = 32'b00000010101101011100111000001100;
   assign mem[1630] = 32'b00000011111110010010001111110100;
   assign mem[1631] = 32'b00001011111101001000100101110000;
   assign mem[1632] = 32'b11111000100010011100110110100000;
   assign mem[1633] = 32'b11110010110100111001100111100000;
   assign mem[1634] = 32'b00000001100001100100001100100100;
   assign mem[1635] = 32'b11111111111110101011101010010110;
   assign mem[1636] = 32'b00001111010111110111101001110000;
   assign mem[1637] = 32'b11110000111110011011100100010000;
   assign mem[1638] = 32'b11111011111001001001000000101000;
   assign mem[1639] = 32'b11111110101010110000000010011100;
   assign mem[1640] = 32'b00000011000111000011011010000100;
   assign mem[1641] = 32'b11110110011111101110001001000000;
   assign mem[1642] = 32'b00000001101000010110011010001100;
   assign mem[1643] = 32'b00000101101000100000100101011000;
   assign mem[1644] = 32'b11111101111010111001010010110100;
   assign mem[1645] = 32'b11111111100001110011101010001101;
   assign mem[1646] = 32'b11110010110001010010100111100000;
   assign mem[1647] = 32'b00000111011111110011100101101000;
   assign mem[1648] = 32'b00000011001110000000110110001000;
   assign mem[1649] = 32'b00000001011010100011001110011000;
   assign mem[1650] = 32'b00000010001011010100000101010000;
   assign mem[1651] = 32'b11111110110111100111101101000110;
   assign mem[1652] = 32'b11111111011110001010110011100100;
   assign mem[1653] = 32'b00000010001100100100010110000000;
   assign mem[1654] = 32'b00000010100000100111000101011000;
   assign mem[1655] = 32'b11111100000111111101010101101100;
   assign mem[1656] = 32'b11111100010101110010101011000100;
   assign mem[1657] = 32'b11111110100010011111101000101010;
   assign mem[1658] = 32'b11111111101100100111110101011011;
   assign mem[1659] = 32'b11111101001000000001010111111100;
   assign mem[1660] = 32'b11111110011111001111011101100000;
   assign mem[1661] = 32'b00000110000100111111110101110000;
   assign mem[1662] = 32'b00000000101010011000001010001100;
   assign mem[1663] = 32'b00000011110000111011100100010100;
   assign mem[1664] = 32'b11111001001011011000110101111000;
   assign mem[1665] = 32'b00001000010100011010111111000000;
   assign mem[1666] = 32'b11111100001101011001001000110000;
   assign mem[1667] = 32'b00000100110001100000110100110000;
   assign mem[1668] = 32'b11111111011110110100100110111100;
   assign mem[1669] = 32'b11110111100100001101110011010000;
   assign mem[1670] = 32'b11111111110010100010101001110000;
   assign mem[1671] = 32'b11111111001000100111101010011111;
   assign mem[1672] = 32'b11111110000110111101101001011000;
   assign mem[1673] = 32'b00000010001111010001110100001100;
   assign mem[1674] = 32'b11111110111000000100100100101010;
   assign mem[1675] = 32'b11111110100111001101010110100100;
   assign mem[1676] = 32'b11111100010100010010100010111000;
   assign mem[1677] = 32'b11111111000100000000101101111111;
   assign mem[1678] = 32'b00000000101101101011111111000011;
   assign mem[1679] = 32'b00000001100111010111010110011110;
   assign mem[1680] = 32'b11111010100101110111011110111000;
   assign mem[1681] = 32'b11110111010110001001011101110000;
   assign mem[1682] = 32'b00001100011100011100001011000000;
   assign mem[1683] = 32'b00000000000110110001001000010001;
   assign mem[1684] = 32'b11110110110111010110110000100000;
   assign mem[1685] = 32'b00000001111101010111100101100110;
   assign mem[1686] = 32'b11111011011100011011010111101000;
   assign mem[1687] = 32'b11111001011101000000100000111000;
   assign mem[1688] = 32'b11111100000010100011111101011100;
   assign mem[1689] = 32'b11111111011111001100111001101101;
   assign mem[1690] = 32'b11111110101011100011011011011000;
   assign mem[1691] = 32'b00000001001101111110000111111100;
   assign mem[1692] = 32'b11111101011011111101110001110000;
   assign mem[1693] = 32'b00000001110000110100001100010110;
   assign mem[1694] = 32'b11111101000101000111110010101100;
   assign mem[1695] = 32'b00000111001010000010110001110000;
   assign mem[1696] = 32'b00000010011000100111000100110000;
   assign mem[1697] = 32'b11110111111110011001000001000000;
   assign mem[1698] = 32'b00000000011101111010010000100001;
   assign mem[1699] = 32'b11111100000110111011110101110000;
   assign mem[1700] = 32'b11111110011111000010011100001000;
   assign mem[1701] = 32'b11111000111110101011101110100000;
   assign mem[1702] = 32'b00000101100100001001111110111000;
   assign mem[1703] = 32'b00001010010101110000010100000000;
   assign mem[1704] = 32'b11111000000110001100001110110000;
   assign mem[1705] = 32'b11110110011001000101110101110000;
   assign mem[1706] = 32'b11101110011010110010001100000000;
   assign mem[1707] = 32'b00010000101011011101001110100000;
   assign mem[1708] = 32'b00000110100001011110101000010000;
   assign mem[1709] = 32'b11101100000011110110010011000000;
   assign mem[1710] = 32'b11111111001011010001011000001001;
   assign mem[1711] = 32'b00001011000100001010110000100000;
   assign mem[1712] = 32'b11111111001011100101010000011010;
   assign mem[1713] = 32'b00000000000110111001101010001001;
   assign mem[1714] = 32'b00001100000100000001011100100000;
   assign mem[1715] = 32'b11111010011110001010110100111000;
   assign mem[1716] = 32'b00000011111010111110001100110100;
   assign mem[1717] = 32'b00000000011011111111010001111001;
   assign mem[1718] = 32'b11111100001000110000001001011100;
   assign mem[1719] = 32'b11101010100001100001111001100000;
   assign mem[1720] = 32'b11111110111000111001011110100010;
   assign mem[1721] = 32'b00000011010110100110111010110000;
   assign mem[1722] = 32'b11110101010101000101001000110000;
   assign mem[1723] = 32'b00000000101001001111001110001010;
   assign mem[1724] = 32'b11111100101111100011000100010100;
   assign mem[1725] = 32'b00001010101001111000001000110000;
   assign mem[1726] = 32'b11111010111000111000110100111000;
   assign mem[1727] = 32'b11111111110100111010001100110000;
   assign mem[1728] = 32'b00000111000100011000100110001000;
   assign mem[1729] = 32'b11111010111000001100111000101000;
   assign mem[1730] = 32'b11111101110110100101101100001000;
   assign mem[1731] = 32'b00000000001111000110011100101101;
   assign mem[1732] = 32'b00000101001110010110110000111000;
   assign mem[1733] = 32'b00000100000111100101001011110000;
   assign mem[1734] = 32'b00000100011100111001111110111000;
   assign mem[1735] = 32'b11110000110010111000110101000000;
   assign mem[1736] = 32'b11111111000001100100100111111000;
   assign mem[1737] = 32'b11111001111110110101000010110000;
   assign mem[1738] = 32'b00000000000101011010101111111110;
   assign mem[1739] = 32'b00000100101110111110111000100000;
   assign mem[1740] = 32'b11110010111011100110111010100000;
   assign mem[1741] = 32'b00000011000110010001110001001100;
   assign mem[1742] = 32'b00001010010100101000000111110000;
   assign mem[1743] = 32'b00000001011110011000010001101110;
   assign mem[1744] = 32'b00000111001110000100000111101000;
   assign mem[1745] = 32'b11111011111010100111011001111000;
   assign mem[1746] = 32'b11111110101110011001110010100100;
   assign mem[1747] = 32'b11100000101001011001010001000000;
   assign mem[1748] = 32'b00000001100111010011100111100110;
   assign mem[1749] = 32'b11100110000001101010000001100000;
   assign mem[1750] = 32'b11111100011111110111001010101000;
   assign mem[1751] = 32'b11111100011110010010010110010000;
   assign mem[1752] = 32'b00000001111110010011100111111010;
   assign mem[1753] = 32'b11111101100000001101101101110100;
   assign mem[1754] = 32'b11111111110001100001101001111000;
   assign mem[1755] = 32'b11111101001101010001110110000100;
   assign mem[1756] = 32'b11111110110101100100111001111010;
   assign mem[1757] = 32'b00000010110001010000111000000100;
   assign mem[1758] = 32'b00000000010101110111011010110101;
   assign mem[1759] = 32'b11111101010010010000100110010000;
   assign mem[1760] = 32'b00000110110010000101111110110000;
   assign mem[1761] = 32'b11111001001000111011001010100000;
   assign mem[1762] = 32'b00000111100111110000100110110000;
   assign mem[1763] = 32'b11111011011100001111011100110000;
   assign mem[1764] = 32'b11110010101001010110000100010000;
   assign mem[1765] = 32'b00000111001010001100110010011000;
   assign mem[1766] = 32'b11111000011010001011010000001000;
   assign mem[1767] = 32'b00000000100000010110000111001100;
   assign mem[1768] = 32'b00000000001010100000011001000110;
   assign mem[1769] = 32'b00000010001010001100011001010100;
   assign mem[1770] = 32'b11111111100110011001111001011110;
   assign mem[1771] = 32'b11111110110110111101010101011110;
   assign mem[1772] = 32'b11111111110101011001101110001111;
   assign mem[1773] = 32'b11111001110011010000000110110000;
   assign mem[1774] = 32'b11111110111100101000010001100110;
   assign mem[1775] = 32'b11111110001010100111000010100100;
   assign mem[1776] = 32'b11111101111111000000111001010100;
   assign mem[1777] = 32'b11111100000110011111101000011000;
   assign mem[1778] = 32'b00000000001011000001000100000100;
   assign mem[1779] = 32'b00000000111011011101010101111011;
   assign mem[1780] = 32'b00000000011100110001010000100111;
   assign mem[1781] = 32'b00000101001001101000010011000000;
   assign mem[1782] = 32'b00000110101000011010100011111000;
   assign mem[1783] = 32'b11111111010111101011010101001001;
   assign mem[1784] = 32'b11111110001100010011111111010110;
   assign mem[1785] = 32'b11111101110101110110011011000100;
   assign mem[1786] = 32'b11111111101110110100001010010011;
   assign mem[1787] = 32'b11110110101000000110001001100000;
   assign mem[1788] = 32'b00000000111010101101011101111010;
   assign mem[1789] = 32'b00000001010010111100010101101100;
   assign mem[1790] = 32'b00000010111100001001010101100100;
   assign mem[1791] = 32'b00000110001010010001100100011000;
   assign mem[1792] = 32'b11111100100110001011000111001000;
   assign mem[1793] = 32'b00000101010001000001011001111000;
   assign mem[1794] = 32'b00000001111111011100001000001100;
   assign mem[1795] = 32'b11111101011101110000101001111000;
   assign mem[1796] = 32'b00000010011010110101000011111000;
   assign mem[1797] = 32'b11110010101001011101111001000000;
   assign mem[1798] = 32'b11111110000010000100101110000100;
   assign mem[1799] = 32'b11111001000111001101011111101000;
   assign mem[1800] = 32'b11111110001100000100101101010010;
   assign mem[1801] = 32'b11111010011001000000010101101000;
   assign mem[1802] = 32'b11111110100010001100101010100100;
   assign mem[1803] = 32'b00000111101010110001011101110000;
   assign mem[1804] = 32'b11101110011110111110010011100000;
   assign mem[1805] = 32'b00000100111111110000001011101000;
   assign mem[1806] = 32'b00000000001100101100101100001111;
   assign mem[1807] = 32'b00000100110000011111011101000000;
   assign mem[1808] = 32'b00000000101000011000111000000010;
   assign mem[1809] = 32'b00000001000001110000110001111000;
   assign mem[1810] = 32'b11111101000000100101010111001100;
   assign mem[1811] = 32'b11110111100001011001110111010000;
   assign mem[1812] = 32'b00000000010001001111100100000110;
   assign mem[1813] = 32'b00000100110010000001101101010000;
   assign mem[1814] = 32'b11110111101101111001101000000000;
   assign mem[1815] = 32'b00000100000101110100111110101000;
   assign mem[1816] = 32'b11110110111000011010110110100000;
   assign mem[1817] = 32'b00000100001111011011111110010000;
   assign mem[1818] = 32'b00000001001110011100111010011110;
   assign mem[1819] = 32'b00000100011010011000001101010000;
   assign mem[1820] = 32'b00000100000010001100001101110000;
   assign mem[1821] = 32'b11111110000110000011000010101110;
   assign mem[1822] = 32'b00000101000001011111000110100000;
   assign mem[1823] = 32'b11111111011111111011011111101101;
   assign mem[1824] = 32'b11100110100010011010001010000000;
   assign mem[1825] = 32'b00000101101111111010001100000000;
   assign mem[1826] = 32'b00000000100101101111111110101001;
   assign mem[1827] = 32'b00000000111101110011010101011010;
   assign mem[1828] = 32'b11111100100110110010100011010100;
   assign mem[1829] = 32'b00000100100101000100110111111000;
   assign mem[1830] = 32'b11111100101111011100111001001000;
   assign mem[1831] = 32'b00001001010100011000010000010000;
   assign mem[1832] = 32'b11110011111101001110000000110000;
   assign mem[1833] = 32'b11110000011100001111010000000000;
   assign mem[1834] = 32'b00010011100001011011011101100000;
   assign mem[1835] = 32'b11111100100111011001001101110000;
   assign mem[1836] = 32'b00001101110011000001100011000000;
   assign mem[1837] = 32'b11100100011011110011001111000000;
   assign mem[1838] = 32'b11111111000101110100000001111001;
   assign mem[1839] = 32'b11101101101010101111001011100000;
   assign mem[1840] = 32'b11111010101101101011100111000000;
   assign mem[1841] = 32'b00000101100001000010111111110000;
   assign mem[1842] = 32'b11111111001100000101010100010000;
   assign mem[1843] = 32'b00001011000011010110100001100000;
   assign mem[1844] = 32'b11111101110111011000011011101000;
   assign mem[1845] = 32'b11111000111000000011011110011000;
   assign mem[1846] = 32'b00001000100011010111010010110000;
   assign mem[1847] = 32'b11110001101101010011100100100000;
   assign mem[1848] = 32'b00000100101000101011001110010000;
   assign mem[1849] = 32'b11110000101101000000010110110000;
   assign mem[1850] = 32'b11111000010011011100101001001000;
   assign mem[1851] = 32'b00000001010001001110001111011010;
   assign mem[1852] = 32'b00000011100100111110111101110100;
   assign mem[1853] = 32'b00001010100010001100101010000000;
   assign mem[1854] = 32'b00000000111110100110000001001100;
   assign mem[1855] = 32'b11110101111100100001001011000000;
   assign mem[1856] = 32'b11111100001101001110110111001100;
   assign mem[1857] = 32'b11111111010011100100100101101010;
   assign mem[1858] = 32'b00000011111100001110010010000000;
   assign mem[1859] = 32'b11101000011011010100110111000000;
   assign mem[1860] = 32'b00000011110000101001100010011100;
   assign mem[1861] = 32'b00000100000011100000111110100000;
   assign mem[1862] = 32'b11111111011000101010000010101110;
   assign mem[1863] = 32'b00000000110000011011010010101111;
   assign mem[1864] = 32'b00000010011111100111111100111000;
   assign mem[1865] = 32'b11111111011011000111001101110110;
   assign mem[1866] = 32'b11111110010001111101001110101000;
   assign mem[1867] = 32'b00000000101101001000100010001000;
   assign mem[1868] = 32'b11111100101010001110110100000000;
   assign mem[1869] = 32'b00000000001010110011001001110010;
   assign mem[1870] = 32'b00000010000011110101000001011000;
   assign mem[1871] = 32'b00000100011100000111010101110000;
   assign mem[1872] = 32'b00000101000100111011101011000000;
   assign mem[1873] = 32'b00000011000001111101111011100000;
   assign mem[1874] = 32'b00000000000110100101011100111000;
   assign mem[1875] = 32'b11111101010010101010010101110100;
   assign mem[1876] = 32'b11111100000010111011011011100000;
   assign mem[1877] = 32'b00000000100100001000100010100110;
   assign mem[1878] = 32'b00000000101111100111001101011000;
   assign mem[1879] = 32'b00000011110100110110111000010000;
   assign mem[1880] = 32'b11111111110111001011111011010000;
   assign mem[1881] = 32'b00000001111001101001001100011110;
   assign mem[1882] = 32'b00000000111101000011001100001001;
   assign mem[1883] = 32'b11111110000010110001100101111000;
   assign mem[1884] = 32'b00000000101010011101001101100101;
   assign mem[1885] = 32'b11111110111011111001110000001000;
   assign mem[1886] = 32'b11111010101000011101111000001000;
   assign mem[1887] = 32'b00000010010110011101100111000000;
   assign mem[1888] = 32'b00000010000010010010111110100100;
   assign mem[1889] = 32'b00000010111000001001100010110000;
   assign mem[1890] = 32'b11111101100000000000100100110000;
   assign mem[1891] = 32'b00000000011111100110001010110111;
   assign mem[1892] = 32'b00000001100111001110101011000100;
   assign mem[1893] = 32'b11111000110011111101100001110000;
   assign mem[1894] = 32'b00000000011001000010011111001111;
   assign mem[1895] = 32'b11111110011101100000001000010110;
   assign mem[1896] = 32'b00000100100100011011110100000000;
   assign mem[1897] = 32'b11111001001111101101111010110000;
   assign mem[1898] = 32'b00000000000101000100010010110111;
   assign mem[1899] = 32'b00000011100111100101001110011000;
   assign mem[1900] = 32'b00000000010100111000010101011100;
   assign mem[1901] = 32'b00000110010011000010011001110000;
   assign mem[1902] = 32'b11111100101001010011010001010000;
   assign mem[1903] = 32'b11111010111001110011100011000000;
   assign mem[1904] = 32'b00000100100001001101000001100000;
   assign mem[1905] = 32'b00000011100001100000000001100100;
   assign mem[1906] = 32'b00000110100101101001101110110000;
   assign mem[1907] = 32'b11110011011100011111111010000000;
   assign mem[1908] = 32'b11111001101100110101100000000000;
   assign mem[1909] = 32'b11111111000011000110111111011010;
   assign mem[1910] = 32'b00000000100101100111011110011100;
   assign mem[1911] = 32'b00000111011010100010110101111000;
   assign mem[1912] = 32'b11111001100110100101000110001000;
   assign mem[1913] = 32'b11111010101011110111100101001000;
   assign mem[1914] = 32'b00001000001000111011001100000000;
   assign mem[1915] = 32'b00000110001000100011011000101000;
   assign mem[1916] = 32'b00000010111101101011000010100100;
   assign mem[1917] = 32'b00000000101101000000111101011111;
   assign mem[1918] = 32'b11111010111111101001100010110000;
   assign mem[1919] = 32'b11110111001110101101100000110000;
   assign mem[1920] = 32'b11111111100100101001100100000000;
   assign mem[1921] = 32'b11111010101011101000111001001000;
   assign mem[1922] = 32'b11111110011011010111111101101010;
   assign mem[1923] = 32'b00000110011111111100001011011000;
   assign mem[1924] = 32'b11111110000100000001101100100010;
   assign mem[1925] = 32'b11111111100110011001110110000010;
   assign mem[1926] = 32'b11111010010101101101110011001000;
   assign mem[1927] = 32'b00000011011101001010010010101000;
   assign mem[1928] = 32'b00000001001100010111001000101100;
   assign mem[1929] = 32'b00000001110010100110110000101100;
   assign mem[1930] = 32'b00000001011011000101010001010110;
   assign mem[1931] = 32'b00000000101100001110110100111010;
   assign mem[1932] = 32'b00000001001110111000001001011010;
   assign mem[1933] = 32'b00000001101110100111001010111100;
   assign mem[1934] = 32'b00000100011101111001111111101000;
   assign mem[1935] = 32'b11111010010010110100111101100000;
   assign mem[1936] = 32'b11111010011011011101101100000000;
   assign mem[1937] = 32'b11111101110100000111011000000100;
   assign mem[1938] = 32'b00000001010101000011110011000000;
   assign mem[1939] = 32'b00000000010010100110110000010111;
   assign mem[1940] = 32'b00000101111100001101000011010000;
   assign mem[1941] = 32'b11110100011100000110000110010000;
   assign mem[1942] = 32'b00000100101110010111111100100000;
   assign mem[1943] = 32'b00000101100010011100010101000000;
   assign mem[1944] = 32'b11110010011011011000101110100000;
   assign mem[1945] = 32'b11111110110100010110001100101010;
   assign mem[1946] = 32'b11111110101011011000010110101110;
   assign mem[1947] = 32'b00000001000011111111001011001110;
   assign mem[1948] = 32'b00000010000110110101111000001000;
   assign mem[1949] = 32'b00000001010010111101001110110000;
   assign mem[1950] = 32'b11111110111011000101111000110010;
   assign mem[1951] = 32'b00000010011110101011010110010000;
   assign mem[1952] = 32'b11111011110011001101101100101000;
   assign mem[1953] = 32'b00000110000101110101001010101000;
   assign mem[1954] = 32'b11111000111011000110010111100000;
   assign mem[1955] = 32'b00000001101011001110101011000000;
   assign mem[1956] = 32'b11111011100110111101101011110000;
   assign mem[1957] = 32'b11111011000010100101010001000000;
   assign mem[1958] = 32'b11111010110001011110001011011000;
   assign mem[1959] = 32'b11111110111010100011000110100000;
   assign mem[1960] = 32'b11111101110001000000000000000100;
   assign mem[1961] = 32'b00001001111001111101100100100000;
   assign mem[1962] = 32'b11111001110001111010111111000000;
   assign mem[1963] = 32'b11110011110011010010101111000000;
   assign mem[1964] = 32'b11111010111100011011111111000000;
   assign mem[1965] = 32'b00001110000111111110011011100000;
   assign mem[1966] = 32'b00000110010110111011110001011000;
   assign mem[1967] = 32'b11111110001101101111001100110110;
   assign mem[1968] = 32'b11111010101010000100011001101000;
   assign mem[1969] = 32'b11100110111100000001011111000000;
   assign mem[1970] = 32'b00000000000010010010101001100111;
   assign mem[1971] = 32'b00000011000010111011101101101100;
   assign mem[1972] = 32'b00000001010001100100001000101110;
   assign mem[1973] = 32'b11110111111010011111011000010000;
   assign mem[1974] = 32'b11111000111001101100011000010000;
   assign mem[1975] = 32'b11111101010101110010101011110100;
   assign mem[1976] = 32'b00000100010101111101001001101000;
   assign mem[1977] = 32'b11111001011110100101010100001000;
   assign mem[1978] = 32'b00000010100000000101011100010000;
   assign mem[1979] = 32'b11111001111000111001100110101000;
   assign mem[1980] = 32'b11110111001000100010010001110000;
   assign mem[1981] = 32'b00001010110110011101000011000000;
   assign mem[1982] = 32'b11110100100000101011110000100000;
   assign mem[1983] = 32'b00000100111111010011100011000000;
   assign mem[1984] = 32'b00000101000100100101101000110000;
   assign mem[1985] = 32'b11111001100111101010111100010000;
   assign mem[1986] = 32'b00000110011010010111111101011000;
   assign mem[1987] = 32'b11111011101111110010110001110000;
   assign mem[1988] = 32'b11111001001010100101111001001000;
   assign mem[1989] = 32'b11110001011000100101100001110000;
   assign mem[1990] = 32'b11110110110001001010111011110000;
   assign mem[1991] = 32'b00001000000111101011110000010000;
   assign mem[1992] = 32'b11110001100010101011101100100000;
   assign mem[1993] = 32'b11110010111010111101110000100000;
   assign mem[1994] = 32'b00000111110100111010001101111000;
   assign mem[1995] = 32'b11111111111111000101101101000100;
   assign mem[1996] = 32'b00000101101001100101110001001000;
   assign mem[1997] = 32'b00000000001101011010000100110000;
   assign mem[1998] = 32'b11111111110000010101111111111100;
   assign mem[1999] = 32'b11110110101001000111111010010000;
   assign mem[2000] = 32'b00000001100001110111010100000010;
   assign mem[2001] = 32'b00000010000000000011000101010000;
   assign mem[2002] = 32'b11111111010111000100101110111101;
   assign mem[2003] = 32'b00000001010011101111011101000000;
   assign mem[2004] = 32'b00000001001010100111100010000010;
   assign mem[2005] = 32'b11111110011010100100000011010000;
   assign mem[2006] = 32'b11111011010001100000001010011000;
   assign mem[2007] = 32'b00000001010100111010001110111100;
   assign mem[2008] = 32'b00000001101010000111100000101010;
   assign mem[2009] = 32'b00000001111110011101100001010100;
   assign mem[2010] = 32'b11111011101111011011001001110000;
   assign mem[2011] = 32'b00010001111111001010011111100000;
   assign mem[2012] = 32'b11110010001111010011111111110000;
   assign mem[2013] = 32'b11111011010001101011000110011000;
   assign mem[2014] = 32'b00001010110110100010101011110000;
   assign mem[2015] = 32'b00000000101010010011000010000111;
   assign mem[2016] = 32'b00000010100100110000011111000100;
   assign mem[2017] = 32'b11101101001100110010000100000000;
   assign mem[2018] = 32'b11111111110111100110111011001101;
   assign mem[2019] = 32'b11110011000001101001011101100000;
   assign mem[2020] = 32'b11111010101001101011010010011000;
   assign mem[2021] = 32'b11111100001101011111110111110000;
   assign mem[2022] = 32'b00000010111000000001101111011100;
   assign mem[2023] = 32'b11111110111101001100111010011100;
   assign mem[2024] = 32'b11110111001010110100101110100000;
   assign mem[2025] = 32'b00000010110010111111110111110100;
   assign mem[2026] = 32'b11111101101110111111100101100000;
   assign mem[2027] = 32'b11111111110010000111101111101000;
   assign mem[2028] = 32'b00000001001100110001100001000000;
   assign mem[2029] = 32'b00000010111001011010101111101100;
   assign mem[2030] = 32'b11111101000100000100100101010000;
   assign mem[2031] = 32'b11111001010110100111011001110000;
   assign mem[2032] = 32'b11111111111011001010101101100001;
   assign mem[2033] = 32'b00000001010001111101001011111100;
   assign mem[2034] = 32'b00000001001100110100000111100100;
   assign mem[2035] = 32'b11111011100101101000100010101000;
   assign mem[2036] = 32'b11111110100100110011011011111100;
   assign mem[2037] = 32'b11111111011101011000000100011010;
   assign mem[2038] = 32'b11111111000010011110011000010101;
   assign mem[2039] = 32'b00000010001111111001011011110000;
   assign mem[2040] = 32'b11111011110101010101110001011000;
   assign mem[2041] = 32'b11111011100011000011010101001000;
   assign mem[2042] = 32'b00000000001001110111001100000110;
   assign mem[2043] = 32'b00000110000000010000010111000000;
   assign mem[2044] = 32'b11111000101111110010001010010000;
   assign mem[2045] = 32'b00000011100011110001110101101100;
   assign mem[2046] = 32'b11111001010101000110011101010000;
   assign mem[2047] = 32'b00000010110001000110111101001000;
   assign mem[2048] = 32'b00000000011110111100100110101111;
   assign mem[2049] = 32'b00000011100100011100000111100000;
   assign mem[2050] = 32'b11111101100000011101100010100100;
   assign mem[2051] = 32'b11111110001000011001000001010110;
   assign mem[2052] = 32'b11111110101101100100000101000110;
   assign mem[2053] = 32'b00000001100001001100000000011000;
   assign mem[2054] = 32'b11111101001010111001110100001000;
   assign mem[2055] = 32'b00000010011011110000110000000100;
   assign mem[2056] = 32'b11111101011111110110100001010000;
   assign mem[2057] = 32'b00000000111000010001010110101111;
   assign mem[2058] = 32'b00000000001011000001000111011111;
   assign mem[2059] = 32'b00000100010100001101101100010000;
   assign mem[2060] = 32'b00000011010000001111101010010100;
   assign mem[2061] = 32'b11111101110100100100100100011100;
   assign mem[2062] = 32'b11111101110010000011010000101000;
   assign mem[2063] = 32'b00000011011000100000000111010100;
   assign mem[2064] = 32'b11101110100101011111000101100000;
   assign mem[2065] = 32'b00000000100011110011111110011000;
   assign mem[2066] = 32'b11111101011000010010011000011000;
   assign mem[2067] = 32'b00000111000110001100110110000000;
   assign mem[2068] = 32'b11111100101100101110000111000100;
   assign mem[2069] = 32'b00000010100000110011011111011000;
   assign mem[2070] = 32'b11111101000111100001101111001100;
   assign mem[2071] = 32'b00000101000010001110101110100000;
   assign mem[2072] = 32'b11111010111100010010110001110000;
   assign mem[2073] = 32'b11101101011101100011100010000000;
   assign mem[2074] = 32'b00001001101000000110101100010000;
   assign mem[2075] = 32'b11111111111011110010111100000110;
   assign mem[2076] = 32'b00000101111010101101101011101000;
   assign mem[2077] = 32'b11110111101001110010111001000000;
   assign mem[2078] = 32'b00000010010000111001010011010000;
   assign mem[2079] = 32'b11111000110101100000010100111000;
   assign mem[2080] = 32'b11111101111110011100000010000100;
   assign mem[2081] = 32'b00000000110010111110100000000001;
   assign mem[2082] = 32'b11111100110011111000001101100100;
   assign mem[2083] = 32'b11111101111011110111011001101000;
   assign mem[2084] = 32'b11111010101010100001000111010000;
   assign mem[2085] = 32'b00001011001010110001011100010000;
   assign mem[2086] = 32'b11111100011111010100011100000000;
   assign mem[2087] = 32'b11111101000100010111010100111100;
   assign mem[2088] = 32'b11111100100101100111111110101000;
   assign mem[2089] = 32'b11111101101000010110111101010100;
   assign mem[2090] = 32'b00000000101110101111011011000010;
   assign mem[2091] = 32'b11111011110010100110110011011000;
   assign mem[2092] = 32'b00000011011111101001110011011100;
   assign mem[2093] = 32'b00000110110011011000001001010000;
   assign mem[2094] = 32'b11101001111100100001110010000000;
   assign mem[2095] = 32'b11111111011011110110000111110101;
   assign mem[2096] = 32'b11111101111011001010000110110100;
   assign mem[2097] = 32'b11111110111100100111011010100100;
   assign mem[2098] = 32'b00000010101000110001011100011000;
   assign mem[2099] = 32'b00000000111011010110000010110000;
   assign mem[2100] = 32'b00000000111001110111001001001101;
   assign mem[2101] = 32'b00000001100101101110111100101010;
   assign mem[2102] = 32'b00000011101010111011000111110000;
   assign mem[2103] = 32'b11111111010011000001000100011111;
   assign mem[2104] = 32'b00000000010100011000100101101100;
   assign mem[2105] = 32'b11110110101011001101111000000000;
   assign mem[2106] = 32'b11111011001100101000011001000000;
   assign mem[2107] = 32'b11111111101010001110101101010000;
   assign mem[2108] = 32'b11111010011000101111110001110000;
   assign mem[2109] = 32'b00000010101100011100100011110000;
   assign mem[2110] = 32'b11111111100101001001010110101001;
   assign mem[2111] = 32'b11111101111100001101110111111100;
   assign mem[2112] = 32'b00000011100000110101100111100100;
   assign mem[2113] = 32'b11111111011110010111001111001001;
   assign mem[2114] = 32'b11111100000010111000111101111100;
   assign mem[2115] = 32'b00000010011000101000101011010000;
   assign mem[2116] = 32'b11111011010011111100110101010000;
   assign mem[2117] = 32'b00000000111100110100010010111001;
   assign mem[2118] = 32'b11111110111011111110000100011110;
   assign mem[2119] = 32'b00000100110011001110011001011000;
   assign mem[2120] = 32'b11111101010000101011111011001000;
   assign mem[2121] = 32'b00000001010011101011101001011100;
   assign mem[2122] = 32'b00000010110001110110011000001000;
   assign mem[2123] = 32'b11111011011010001001000010110000;
   assign mem[2124] = 32'b00000111010100110111101110101000;
   assign mem[2125] = 32'b00000000101101111101101110101000;
   assign mem[2126] = 32'b00000001111011001111001010001000;
   assign mem[2127] = 32'b11110100001111010000001111000000;
   assign mem[2128] = 32'b00000010011100100101100100011100;
   assign mem[2129] = 32'b11110001110100100001100111000000;
   assign mem[2130] = 32'b00000000001100111010110101011111;
   assign mem[2131] = 32'b11111111101101011111001101000111;
   assign mem[2132] = 32'b00000000010001001011001010100010;
   assign mem[2133] = 32'b11111100011111011010010110101100;
   assign mem[2134] = 32'b11111010110000000001011010101000;
   assign mem[2135] = 32'b00000100000010001010100100101000;
   assign mem[2136] = 32'b00000000100001100101011100010011;
   assign mem[2137] = 32'b00000011001010011010010000110100;
   assign mem[2138] = 32'b11111111010011110100110111111011;
   assign mem[2139] = 32'b00000011000101100010101000011100;
   assign mem[2140] = 32'b11111101000100101110000110010100;
   assign mem[2141] = 32'b00000011000100010001000101011100;
   assign mem[2142] = 32'b11110110000001111010100010000000;
   assign mem[2143] = 32'b11111001100111100100000011100000;
   assign mem[2144] = 32'b00001000101111101011010111010000;
   assign mem[2145] = 32'b11111011110000111100110100111000;
   assign mem[2146] = 32'b00000111011010000110001111000000;
   assign mem[2147] = 32'b00000110000000001000111111101000;
   assign mem[2148] = 32'b11111101111111101000011110100000;
   assign mem[2149] = 32'b11111001000001001011110010001000;
   assign mem[2150] = 32'b00000111100110010110111000001000;
   assign mem[2151] = 32'b11111101000111000011001100010000;
   assign mem[2152] = 32'b00000111111101010011011100010000;
   assign mem[2153] = 32'b00000010000000101101010010110000;
   assign mem[2154] = 32'b00000110111100101111010110101000;
   assign mem[2155] = 32'b11110111100000001101100010100000;
   assign mem[2156] = 32'b11111010000001001010111011011000;
   assign mem[2157] = 32'b11111111001101000011011000010011;
   assign mem[2158] = 32'b11111100010001011111001100100100;
   assign mem[2159] = 32'b11111100001110001111100100110100;
   assign mem[2160] = 32'b00000100011111100111101000110000;
   assign mem[2161] = 32'b00000001100101111100001001111000;
   assign mem[2162] = 32'b00000100011111101100111011010000;
   assign mem[2163] = 32'b00000010111010000100010001001000;
   assign mem[2164] = 32'b00001100110000100101100011100000;
   assign mem[2165] = 32'b11110111110101111100101111010000;
   assign mem[2166] = 32'b11111110000001110101011111111010;
   assign mem[2167] = 32'b11111000011111110110100101000000;
   assign mem[2168] = 32'b00000010101011010011100010011100;
   assign mem[2169] = 32'b11110000011010100000010010000000;
   assign mem[2170] = 32'b11111101110111010010110001001000;
   assign mem[2171] = 32'b00000111100001001011100000000000;
   assign mem[2172] = 32'b00000110100111100001001110110000;
   assign mem[2173] = 32'b00000110001000100111001010011000;
   assign mem[2174] = 32'b11111101001101110111100101101000;
   assign mem[2175] = 32'b11110001101100101001000111010000;
   assign mem[2176] = 32'b00000100000011010001100111101000;
   assign mem[2177] = 32'b11111101001100100111100110101000;
   assign mem[2178] = 32'b11111010001011110010001011100000;
   assign mem[2179] = 32'b11110111001110011001001010010000;
   assign mem[2180] = 32'b11111001010111011010000011000000;
   assign mem[2181] = 32'b00001000011001101110111010010000;
   assign mem[2182] = 32'b00000010110101000101010010111000;
   assign mem[2183] = 32'b11111000011110100100001001110000;
   assign mem[2184] = 32'b00000101101111000110000101111000;
   assign mem[2185] = 32'b11111000010101111010100000111000;
   assign mem[2186] = 32'b11111110101101010101000000100000;
   assign mem[2187] = 32'b11111100000000101011010011001000;
   assign mem[2188] = 32'b11111110110010110000110010110110;
   assign mem[2189] = 32'b11110101111001100110010111100000;
   assign mem[2190] = 32'b00000011001101001000101111100000;
   assign mem[2191] = 32'b00000100111001000001001110110000;
   assign mem[2192] = 32'b11111011011101111111000100101000;
   assign mem[2193] = 32'b11110111111101100010011100010000;
   assign mem[2194] = 32'b00000101111011111001101000011000;
   assign mem[2195] = 32'b00000100100010101101101110111000;
   assign mem[2196] = 32'b00000000110100110000000010001101;
   assign mem[2197] = 32'b11111100100111101110101010100100;
   assign mem[2198] = 32'b00000001111100100110010100100010;
   assign mem[2199] = 32'b00000000100110010100101010000010;
   assign mem[2200] = 32'b11111101110100011001010010010000;
   assign mem[2201] = 32'b11111110001110100011001111010010;
   assign mem[2202] = 32'b11111101101101000110100000010000;
   assign mem[2203] = 32'b00000000111001100001010111001001;
   assign mem[2204] = 32'b11110101011011001001000100100000;
   assign mem[2205] = 32'b00000001110110010001100001000110;
   assign mem[2206] = 32'b11111010000000010100011110001000;
   assign mem[2207] = 32'b00000101001110101001001010110000;
   assign mem[2208] = 32'b00000000001100110010110011001100;
   assign mem[2209] = 32'b00000001110110010101101000111100;
   assign mem[2210] = 32'b11111110011010010100000111011000;
   assign mem[2211] = 32'b11111011010101010111011001010000;
   assign mem[2212] = 32'b11111101010011101110001110001100;
   assign mem[2213] = 32'b00000000100000101010110110010001;
   assign mem[2214] = 32'b11111001100110000000100000101000;
   assign mem[2215] = 32'b11111110111110001000010111011100;
   assign mem[2216] = 32'b11111011000100000110110111010000;
   assign mem[2217] = 32'b00000011000010110000000001101000;
   assign mem[2218] = 32'b00000000011100000111111110000101;
   assign mem[2219] = 32'b00000001011111111110111111101110;
   assign mem[2220] = 32'b11111101011101110000001010101000;
   assign mem[2221] = 32'b00000101001001011101011010001000;
   assign mem[2222] = 32'b00000110011111010000111000001000;
   assign mem[2223] = 32'b11111111010001110001101100000111;
   assign mem[2224] = 32'b00001010001000110100111110110000;
   assign mem[2225] = 32'b11111101001011100111000001011100;
   assign mem[2226] = 32'b00000010101111100110011101101000;
   assign mem[2227] = 32'b00000000000110111011001110010011;
   assign mem[2228] = 32'b11111000101010000000111111110000;
   assign mem[2229] = 32'b11110101111101010010111100010000;
   assign mem[2230] = 32'b11111110101111101010101101001110;
   assign mem[2231] = 32'b11111010011001111001110011011000;
   assign mem[2232] = 32'b11111110110110101101101101011010;
   assign mem[2233] = 32'b11111101110100001110010110010100;
   assign mem[2234] = 32'b11110010010011101111011101110000;
   assign mem[2235] = 32'b00000110111111110111101110111000;
   assign mem[2236] = 32'b00000011011011000100100110011100;
   assign mem[2237] = 32'b00000001001000100001110011010110;
   assign mem[2238] = 32'b11111100011101101000010010101000;
   assign mem[2239] = 32'b00000101100010010010111010010000;
   assign mem[2240] = 32'b00000000100001110000101100010001;
   assign mem[2241] = 32'b00001000111110000111001101100000;
   assign mem[2242] = 32'b11111111000111001111110101001010;
   assign mem[2243] = 32'b00000000110001101101001111101010;
   assign mem[2244] = 32'b11111110000010111011111010000110;
   assign mem[2245] = 32'b00000000010000000001110000100101;
   assign mem[2246] = 32'b00000001111010000100100110011010;
   assign mem[2247] = 32'b00000001010101100001100110000100;
   assign mem[2248] = 32'b11111011100000001110010000011000;
   assign mem[2249] = 32'b00000000101111110100110111111010;
   assign mem[2250] = 32'b00001000001100111111001110110000;
   assign mem[2251] = 32'b00000111111101111101010001100000;
   assign mem[2252] = 32'b11110101110101101011000011110000;
   assign mem[2253] = 32'b11110011101011011010101000110000;
   assign mem[2254] = 32'b00000111000100011100101101111000;
   assign mem[2255] = 32'b00000000001000011110010011011111;
   assign mem[2256] = 32'b00000111011100000011110111000000;
   assign mem[2257] = 32'b11111101111110110011010111001100;
   assign mem[2258] = 32'b00000000101001101000100001000001;
   assign mem[2259] = 32'b11111011000000011011111101010000;
   assign mem[2260] = 32'b11111001011101101110110101000000;
   assign mem[2261] = 32'b11110000101111110101110100010000;
   assign mem[2262] = 32'b00000000001010010010101000100001;
   assign mem[2263] = 32'b00000010000011101100110111100100;
   assign mem[2264] = 32'b11101000011111101000000000000000;
   assign mem[2265] = 32'b00000110011001010011111001111000;
   assign mem[2266] = 32'b00000010110101110111001101011000;
   assign mem[2267] = 32'b11111101011111001100000001101100;
   assign mem[2268] = 32'b00000100110111010101100011100000;
   assign mem[2269] = 32'b00000101000001111110010100101000;
   assign mem[2270] = 32'b11110110110001110001101100000000;
   assign mem[2271] = 32'b00001100010011111010100011110000;
   assign mem[2272] = 32'b11101011000000000010110011000000;
   assign mem[2273] = 32'b00000001101111111111010100000110;
   assign mem[2274] = 32'b00001100110111010011100111010000;
   assign mem[2275] = 32'b11111110100000011011010011101000;
   assign mem[2276] = 32'b00000110111000011001111001111000;
   assign mem[2277] = 32'b11100100111001010011000001000000;
   assign mem[2278] = 32'b00000010111001011010110110000000;
   assign mem[2279] = 32'b11110001011101111101111101110000;
   assign mem[2280] = 32'b11111100111101110011011111100100;
   assign mem[2281] = 32'b00000000101000010000000001101100;
   assign mem[2282] = 32'b11111111011011111111100100100010;
   assign mem[2283] = 32'b00000010100000000100100110101000;
   assign mem[2284] = 32'b11111010111000111111000000110000;
   assign mem[2285] = 32'b11111110000010111101000100100010;
   assign mem[2286] = 32'b11111010100101110010101101111000;
   assign mem[2287] = 32'b11111110001110001010010101110010;
   assign mem[2288] = 32'b00000001010001100001110111111100;
   assign mem[2289] = 32'b00000100001001111111101010101000;
   assign mem[2290] = 32'b11111111000111110110010001100010;
   assign mem[2291] = 32'b11111110001010110000100111010010;
   assign mem[2292] = 32'b00000010100100011101100100111100;
   assign mem[2293] = 32'b00000000110100011110011101011111;
   assign mem[2294] = 32'b11111100001111011000001101001000;
   assign mem[2295] = 32'b11111100110000000111110001101100;
   assign mem[2296] = 32'b11111001101111110101001101010000;
   assign mem[2297] = 32'b00000110001001110001100001011000;
   assign mem[2298] = 32'b00000010101001011101111011010100;
   assign mem[2299] = 32'b00000101010001101010101100110000;
   assign mem[2300] = 32'b11111100011000000101111101000100;
   assign mem[2301] = 32'b00000001100000000101000100101000;
   assign mem[2302] = 32'b11111001011111001000101010001000;
   assign mem[2303] = 32'b11111110000101111110100101011100;
   assign mem[2304] = 32'b00000001010000111111011011001100;
   assign mem[2305] = 32'b00000110101111111111100010111000;
   assign mem[2306] = 32'b11111110111111000010101111101000;
   assign mem[2307] = 32'b00000001001001111100000111111000;
   assign mem[2308] = 32'b00000010001011000101001001010000;
   assign mem[2309] = 32'b11111000011001111010101010101000;
   assign mem[2310] = 32'b11111100111101001101100101100100;
   assign mem[2311] = 32'b00000010011011111000010001100100;
   assign mem[2312] = 32'b11101111001010001101110101100000;
   assign mem[2313] = 32'b11111001101100001100111001111000;
   assign mem[2314] = 32'b00000100100010111001111100110000;
   assign mem[2315] = 32'b00000100111011010101010110110000;
   assign mem[2316] = 32'b11111101011001101001110001010100;
   assign mem[2317] = 32'b00000000011010011101001011000110;
   assign mem[2318] = 32'b11111001000011010011111010000000;
   assign mem[2319] = 32'b00000011100000011101010110001000;
   assign mem[2320] = 32'b00000000000000101000110111000100;
   assign mem[2321] = 32'b11111010110011011010000111001000;
   assign mem[2322] = 32'b00001000010101010011011101000000;
   assign mem[2323] = 32'b00000000111010100000110001010010;
   assign mem[2324] = 32'b11111010100100000011000100010000;
   assign mem[2325] = 32'b11111011010100100011101110100000;
   assign mem[2326] = 32'b11111111100100110011101110011101;
   assign mem[2327] = 32'b11111110110001011000001111000100;
   assign mem[2328] = 32'b11110011100011001110011100110000;
   assign mem[2329] = 32'b00000100110101001100100111100000;
   assign mem[2330] = 32'b11111100000111010101100011011000;
   assign mem[2331] = 32'b00000011010000010110001100100100;
   assign mem[2332] = 32'b11110111100011010001010110000000;
   assign mem[2333] = 32'b11111100101011011110000111001000;
   assign mem[2334] = 32'b11101110010011011001000010100000;
   assign mem[2335] = 32'b00001001000101011110111100110000;
   assign mem[2336] = 32'b00000001001110010100000101100010;
   assign mem[2337] = 32'b11110111100010111101100111100000;
   assign mem[2338] = 32'b00000001100100011010000100100100;
   assign mem[2339] = 32'b00000100110011000101101101000000;
   assign mem[2340] = 32'b11111111000110111100111010011111;
   assign mem[2341] = 32'b11111111111010100011001111000010;
   assign mem[2342] = 32'b11111100010101011100011000010000;
   assign mem[2343] = 32'b00000100100110101111000010000000;
   assign mem[2344] = 32'b11110100011011111000001101010000;
   assign mem[2345] = 32'b00000010111100011001000001011100;
   assign mem[2346] = 32'b11111111001110011001010110000010;
   assign mem[2347] = 32'b00001001001101101001100010110000;
   assign mem[2348] = 32'b11110100100000000101110010000000;
   assign mem[2349] = 32'b11101111101011010100100101000000;
   assign mem[2350] = 32'b11111010101111010000011100010000;
   assign mem[2351] = 32'b00000010100010111110010110010100;
   assign mem[2352] = 32'b00000011101111001111110000100100;
   assign mem[2353] = 32'b00000110011010100100100011100000;
   assign mem[2354] = 32'b00001000001101001001101010000000;
   assign mem[2355] = 32'b11110110111011011001000001000000;
   assign mem[2356] = 32'b11111011111100110001111110101000;
   assign mem[2357] = 32'b00000010100011010001011100100100;
   assign mem[2358] = 32'b00000000000111001011000101111000;
   assign mem[2359] = 32'b11111000100000001000001111111000;
   assign mem[2360] = 32'b11111011000001010101110011101000;
   assign mem[2361] = 32'b00000010001000111010001100100100;
   assign mem[2362] = 32'b11111100000010101001000010000100;
   assign mem[2363] = 32'b00000010001100100001000111110000;
   assign mem[2364] = 32'b00000101101010010110100000100000;
   assign mem[2365] = 32'b00000001001010110011000000111110;
   assign mem[2366] = 32'b11110110111101011010111100110000;
   assign mem[2367] = 32'b00000010000100100101101101110100;
   assign mem[2368] = 32'b00000010000110010001000001010100;
   assign mem[2369] = 32'b11111110011110110111110011011110;
   assign mem[2370] = 32'b00000001100100001001010010011010;
   assign mem[2371] = 32'b11111001011111100011101111111000;
   assign mem[2372] = 32'b00000010110101011111111110111100;
   assign mem[2373] = 32'b00000101010110101001101000010000;
   assign mem[2374] = 32'b11111000111101110010011011100000;
   assign mem[2375] = 32'b11110110011001000000001010000000;
   assign mem[2376] = 32'b11111101010000101010111000100100;
   assign mem[2377] = 32'b00000010100111100011011000011100;
   assign mem[2378] = 32'b00000011100010000100000111000100;
   assign mem[2379] = 32'b00000100011011111000101001001000;
   assign mem[2380] = 32'b11111110010010001100010100010010;
   assign mem[2381] = 32'b00000100101100010001111111011000;
   assign mem[2382] = 32'b00000101011010001000100010101000;
   assign mem[2383] = 32'b00000010000110111111010110101100;
   assign mem[2384] = 32'b00000000010011101100001011100001;
   assign mem[2385] = 32'b00000001110011110100001000011100;
   assign mem[2386] = 32'b11110101111001010001101000010000;
   assign mem[2387] = 32'b11110010011100101001010111000000;
   assign mem[2388] = 32'b11111000001000001110010000000000;
   assign mem[2389] = 32'b11111011010010001010101010000000;
   assign mem[2390] = 32'b11111110110010011001101101100000;
   assign mem[2391] = 32'b00000010100110011001100111011000;
   assign mem[2392] = 32'b11111100111010001100100011111100;
   assign mem[2393] = 32'b11111100101011000000010000000100;
   assign mem[2394] = 32'b00000011000010011100001000110100;
   assign mem[2395] = 32'b11111101001011001000011110011100;
   assign mem[2396] = 32'b00000001101100101010110000110110;
   assign mem[2397] = 32'b00000010011101111111100100001100;
   assign mem[2398] = 32'b11111111110001001010011000010011;
   assign mem[2399] = 32'b11111100001111100101110110000100;
   assign mem[2400] = 32'b00000100001011101000010111100000;
   assign mem[2401] = 32'b11110011110100110110011010010000;
   assign mem[2402] = 32'b11111110010010010011001000101010;
   assign mem[2403] = 32'b00000000101101111111010011011001;
   assign mem[2404] = 32'b11110011111101011111001101000000;
   assign mem[2405] = 32'b00000111001001001010010010100000;
   assign mem[2406] = 32'b00000011100100101001001000111000;
   assign mem[2407] = 32'b11111000101100001111100000011000;
   assign mem[2408] = 32'b00000001111000100011000010100000;
   assign mem[2409] = 32'b11111001110100000010111111100000;
   assign mem[2410] = 32'b11111111101100100100111000011010;
   assign mem[2411] = 32'b00000100010011001011001101111000;
   assign mem[2412] = 32'b11111011111001111001101011111000;
   assign mem[2413] = 32'b11110110011100011100111000110000;
   assign mem[2414] = 32'b00000011101001000011111110100100;
   assign mem[2415] = 32'b00000101010011010011101001001000;
   assign mem[2416] = 32'b00000001001101011000001001001000;
   assign mem[2417] = 32'b11111011010000111111010010000000;
   assign mem[2418] = 32'b11111011010110011111000110000000;
   assign mem[2419] = 32'b00000010101010110001111110110000;
   assign mem[2420] = 32'b11111110100010000111101011101100;
   assign mem[2421] = 32'b00000010110001011110110101111100;
   assign mem[2422] = 32'b00000000001001101100101011000011;
   assign mem[2423] = 32'b11111110100001010011000010000100;
   assign mem[2424] = 32'b00000100011110100001000101101000;
   assign mem[2425] = 32'b00000001010001110100100100000100;
   assign mem[2426] = 32'b00000100100010111101000101110000;
   assign mem[2427] = 32'b11111001101001001100100100110000;
   assign mem[2428] = 32'b11111111110001011000111101000100;
   assign mem[2429] = 32'b11111100111111101100110111000000;
   assign mem[2430] = 32'b00000000000111001110101110101010;
   assign mem[2431] = 32'b00001010110110111110111001010000;
   assign mem[2432] = 32'b11110110111001010100110111010000;
   assign mem[2433] = 32'b11111100101100100111010011011100;
   assign mem[2434] = 32'b00001000100110101001001000110000;
   assign mem[2435] = 32'b11110111100111011111110000000000;
   assign mem[2436] = 32'b00001101011001100000100010000000;
   assign mem[2437] = 32'b11111110000011001011100011010110;
   assign mem[2438] = 32'b00000011110010010100100111001100;
   assign mem[2439] = 32'b11110101111001000100101110010000;
   assign mem[2440] = 32'b00000011101111110111101000000000;
   assign mem[2441] = 32'b11111011111011110010010010000000;
   assign mem[2442] = 32'b11111110000011100011101101100000;
   assign mem[2443] = 32'b00000101010111011111011010000000;
   assign mem[2444] = 32'b11100110011001010010001010100000;
   assign mem[2445] = 32'b00000100100001111111001100000000;
   assign mem[2446] = 32'b00000001111000101011001110101010;
   assign mem[2447] = 32'b11111011111100100011000100111000;
   assign mem[2448] = 32'b00000001010001100100001000011100;
   assign mem[2449] = 32'b00000010111000011101001010111000;
   assign mem[2450] = 32'b00000001001000111001011001001000;
   assign mem[2451] = 32'b11101111110011110100111011000000;
   assign mem[2452] = 32'b11111111111010011000011101110100;
   assign mem[2453] = 32'b00000000010111100010111010100110;
   assign mem[2454] = 32'b11110001000011110110101100100000;
   assign mem[2455] = 32'b00000100010100001010100111000000;
   assign mem[2456] = 32'b11111101001101101001110110101100;
   assign mem[2457] = 32'b00000101001001100110001011010000;
   assign mem[2458] = 32'b00000000010001011000101111010000;
   assign mem[2459] = 32'b00000111011111011000011000001000;
   assign mem[2460] = 32'b11111111001101000000100111010011;
   assign mem[2461] = 32'b11111111101001101010101100000011;
   assign mem[2462] = 32'b11111101011000000110111000000100;
   assign mem[2463] = 32'b11111100011010100000101010101100;
   assign mem[2464] = 32'b11110001100001100000101100100000;
   assign mem[2465] = 32'b00000111010101100010101000001000;
   assign mem[2466] = 32'b00000110100111101001000011111000;
   assign mem[2467] = 32'b11101101010010110011010110100000;
   assign mem[2468] = 32'b11111101011000110100111010110000;
   assign mem[2469] = 32'b00000100001001110100110001100000;
   assign mem[2470] = 32'b11110101100010110001100101010000;
   assign mem[2471] = 32'b00000100010000111000111000010000;
   assign mem[2472] = 32'b11110001110011100011000101010000;
   assign mem[2473] = 32'b00000001100100111010010010011010;
   assign mem[2474] = 32'b00010000001101111000011101100000;
   assign mem[2475] = 32'b00000010100111010100111010000000;
   assign mem[2476] = 32'b00000101101010010111101001001000;
   assign mem[2477] = 32'b11110101100111000111101110000000;
   assign mem[2478] = 32'b00000001000001010101110100101110;
   assign mem[2479] = 32'b11101110100010101010001001100000;
   assign mem[2480] = 32'b11111111110010110001111101110011;
   assign mem[2481] = 32'b00000010011101001101101011000100;
   assign mem[2482] = 32'b00000001110101101100101001011110;
   assign mem[2483] = 32'b00001011110101100100000000010000;
   assign mem[2484] = 32'b11111110001100001100011111001110;
   assign mem[2485] = 32'b11110110110101100010101111110000;
   assign mem[2486] = 32'b11111101001111000110110100110000;
   assign mem[2487] = 32'b00000010111110011100111001000000;
   assign mem[2488] = 32'b11111110000011101101110111001110;
   assign mem[2489] = 32'b11110100011011101001111010010000;
   assign mem[2490] = 32'b00000011000100110110110011110100;
   assign mem[2491] = 32'b11110011011100011110010000100000;
   assign mem[2492] = 32'b00000101001101011011000001110000;
   assign mem[2493] = 32'b00001100001010010001001110110000;
   assign mem[2494] = 32'b11111101111101100111001010100100;
   assign mem[2495] = 32'b11111101101111011111111000110000;
   assign mem[2496] = 32'b11111011010110101101111111011000;
   assign mem[2497] = 32'b11111100011001110000100111100100;
   assign mem[2498] = 32'b11111100111000011111101011010100;
   assign mem[2499] = 32'b11111010111110110011001011011000;
   assign mem[2500] = 32'b00000000000111010101010111100011;
   assign mem[2501] = 32'b00000001100110000100001101110000;
   assign mem[2502] = 32'b11111100111011000111011011111000;
   assign mem[2503] = 32'b00000000001100000101111001100111;
   assign mem[2504] = 32'b11111101010000000010110111101000;
   assign mem[2505] = 32'b11111111011011001011100111111100;
   assign mem[2506] = 32'b11111001001000111111011100100000;
   assign mem[2507] = 32'b11111111001100110111110011010001;
   assign mem[2508] = 32'b11111111011110100011101011011111;
   assign mem[2509] = 32'b11111111111010010110001011100010;
   assign mem[2510] = 32'b00000011010001011101101100100000;
   assign mem[2511] = 32'b11111111011100000100000001111111;
   assign mem[2512] = 32'b00000010001001101110010001110100;
   assign mem[2513] = 32'b11111111011000100011011000011110;
   assign mem[2514] = 32'b11111111010000010100100111101111;
   assign mem[2515] = 32'b11111110111111010101101010101100;
   assign mem[2516] = 32'b11110110100101111011011001100000;
   assign mem[2517] = 32'b11111111001011010110111101111101;
   assign mem[2518] = 32'b00000001001100101011100011011110;
   assign mem[2519] = 32'b00000010010011110111100000001000;
   assign mem[2520] = 32'b00000000110101111011101000110100;
   assign mem[2521] = 32'b00000100100010100101111010001000;
   assign mem[2522] = 32'b00000000010111100010001010010110;
   assign mem[2523] = 32'b11111100110001001100110110100100;
   assign mem[2524] = 32'b00000101000010111000001101001000;
   assign mem[2525] = 32'b00000000001010001000001010010111;
   assign mem[2526] = 32'b11111111011100001110100101001010;
   assign mem[2527] = 32'b11111111100110001100110000101100;
   assign mem[2528] = 32'b00000001010011011011101001100000;
   assign mem[2529] = 32'b00000010011110100011000010011100;
   assign mem[2530] = 32'b00000100010101000101101011010000;
   assign mem[2531] = 32'b00000101010010101000100111010000;
   assign mem[2532] = 32'b11111010100100010011000100110000;
   assign mem[2533] = 32'b11110110000001010101100011110000;
   assign mem[2534] = 32'b00000100010110110000011000111000;
   assign mem[2535] = 32'b11111101011001111100110101001000;
   assign mem[2536] = 32'b00000001001001101101010100010110;
   assign mem[2537] = 32'b00000010110111000101000001111100;
   assign mem[2538] = 32'b11111101000111111010110110110100;
   assign mem[2539] = 32'b00000001000001000110000010110110;
   assign mem[2540] = 32'b11111011111100011100100100101000;
   assign mem[2541] = 32'b00000011011111000101001111110100;
   assign mem[2542] = 32'b00000011010000001110011011100100;
   assign mem[2543] = 32'b11110110001011000001110001110000;
   assign mem[2544] = 32'b00001110101100101100001101010000;
   assign mem[2545] = 32'b11111111000101001101111101110101;
   assign mem[2546] = 32'b00000011001110001111101001110100;
   assign mem[2547] = 32'b11101110110010000111111100000000;
   assign mem[2548] = 32'b00000000010110101111110101111001;
   assign mem[2549] = 32'b11101010001001100100010110100000;
   assign mem[2550] = 32'b11111101111000001111011010100100;
   assign mem[2551] = 32'b00001001011001000001110001000000;
   assign mem[2552] = 32'b11111000010101011001110100110000;
   assign mem[2553] = 32'b00000000011001111010111101001111;
   assign mem[2554] = 32'b00001001110001000111001000100000;
   assign mem[2555] = 32'b00000101010101111100111010011000;
   assign mem[2556] = 32'b00000000101000000110100001010011;
   assign mem[2557] = 32'b11111111000000000100111101010001;
   assign mem[2558] = 32'b11111111001001100000111101001011;
   assign mem[2559] = 32'b11110100011101001110101011000000;
   assign mem[2560] = 32'b00000101000110100000001100111000;
   assign mem[2561] = 32'b11111001101110110100011000111000;
   assign mem[2562] = 32'b11110101011101110110101011110000;
   assign mem[2563] = 32'b11111101000101111110111110011000;
   assign mem[2564] = 32'b11111111010001101011011011011101;
   assign mem[2565] = 32'b11111110111010010010110110011110;
   assign mem[2566] = 32'b11111101111110001001100011011100;
   assign mem[2567] = 32'b00000100101011111011100000010000;
   assign mem[2568] = 32'b00000101101010000110000111101000;
   assign mem[2569] = 32'b00000011011000011010101110100100;
   assign mem[2570] = 32'b11111110110110011010001000001000;
   assign mem[2571] = 32'b00000000101110101011110010010011;
   assign mem[2572] = 32'b11111110101000011110110110110100;
   assign mem[2573] = 32'b00000000011000001100111001010011;
   assign mem[2574] = 32'b00000000000010010010111101011100;
   assign mem[2575] = 32'b11111000001100010111000001011000;
   assign mem[2576] = 32'b11111001100111110111111111111000;
   assign mem[2577] = 32'b11111110011010011001000100010000;
   assign mem[2578] = 32'b00000000101001011110100011101010;
   assign mem[2579] = 32'b00000010000011111010101001110000;
   assign mem[2580] = 32'b00000101100111000110001100100000;
   assign mem[2581] = 32'b11110100101011011011010101000000;
   assign mem[2582] = 32'b00000011000000111001111111101000;
   assign mem[2583] = 32'b00000111110111010100111100011000;
   assign mem[2584] = 32'b11111001110001000110001001001000;
   assign mem[2585] = 32'b11110000101101111110000001110000;
   assign mem[2586] = 32'b00000110011011110000011100100000;
   assign mem[2587] = 32'b00000010111100111101011010010100;
   assign mem[2588] = 32'b00000001111110011010010000011110;
   assign mem[2589] = 32'b00000100001010010001000101100000;
   assign mem[2590] = 32'b11111100101101101100110101101000;
   assign mem[2591] = 32'b11110101001011000010010111010000;
   assign mem[2592] = 32'b11111000010001000111110000001000;
   assign mem[2593] = 32'b11110010100011000001011000010000;
   assign mem[2594] = 32'b11111101110101000111110110011000;
   assign mem[2595] = 32'b00000010101001101010010101010000;
   assign mem[2596] = 32'b11111110011011101110001101100010;
   assign mem[2597] = 32'b11110001111001111100111110010000;
   assign mem[2598] = 32'b00000011000010110001110100010000;
   assign mem[2599] = 32'b11110101011010011011101100000000;
   assign mem[2600] = 32'b11111010011000010010111110000000;
   assign mem[2601] = 32'b00000000010001110110010010000000;
   assign mem[2602] = 32'b11110110001000000001010001010000;
   assign mem[2603] = 32'b11101100010010000011011111000000;
   assign mem[2604] = 32'b11111100101111000001111011111000;
   assign mem[2605] = 32'b00000101001111110000110011011000;
   assign mem[2606] = 32'b00001001101010100001101110010000;
   assign mem[2607] = 32'b11111100011011011010000001001100;
   assign mem[2608] = 32'b11111111011000010001000100110010;
   assign mem[2609] = 32'b11111011001110001111111010101000;
   assign mem[2610] = 32'b00000111111100000101100101001000;
   assign mem[2611] = 32'b00000111111110111010100011111000;
   assign mem[2612] = 32'b11111001011011100001010101111000;
   assign mem[2613] = 32'b11110110111001011000001011110000;
   assign mem[2614] = 32'b00000111110001010111111110000000;
   assign mem[2615] = 32'b00000010000110000100000101011100;
   assign mem[2616] = 32'b00000010111010010101111010101000;
   assign mem[2617] = 32'b11111111110011011000001001010000;
   assign mem[2618] = 32'b11111101101000000000000000010100;
   assign mem[2619] = 32'b11110110110010001110110001010000;
   assign mem[2620] = 32'b11110011110111111000001001010000;
   assign mem[2621] = 32'b11111111100011100100111111111101;
   assign mem[2622] = 32'b11111101011100001110010011000000;
   assign mem[2623] = 32'b00000011010111000101000001001100;
   assign mem[2624] = 32'b11111010100111100100010000100000;
   assign mem[2625] = 32'b00000001010101001111001011110100;
   assign mem[2626] = 32'b00000011011011100100111100011000;
   assign mem[2627] = 32'b00000010011011111001101100100100;
   assign mem[2628] = 32'b00000000111001111110111111111010;
   assign mem[2629] = 32'b11111000010100000000100010111000;
   assign mem[2630] = 32'b11110110111101010011110000110000;
   assign mem[2631] = 32'b00001001111000001010011011100000;
   assign mem[2632] = 32'b11101100011010101010011011100000;
   assign mem[2633] = 32'b11111011111011101111110110000000;
   assign mem[2634] = 32'b00000001001101101010100100001010;
   assign mem[2635] = 32'b00001001010011001001110100010000;
   assign mem[2636] = 32'b00000100010010100101010001110000;
   assign mem[2637] = 32'b00000011001100101101100101001100;
   assign mem[2638] = 32'b11111110011011110101111001000010;
   assign mem[2639] = 32'b00000010000000001110011111100100;
   assign mem[2640] = 32'b11111110101010111111101110111010;
   assign mem[2641] = 32'b00000000010000011001100101010100;
   assign mem[2642] = 32'b11111011111010001110001010100000;
   assign mem[2643] = 32'b11111101111110001001011000010000;
   assign mem[2644] = 32'b11111111111011110011001000111000;
   assign mem[2645] = 32'b11111111001010101010110001101010;
   assign mem[2646] = 32'b11111110010011000101001110001000;
   assign mem[2647] = 32'b00000011001100001101111110000000;
   assign mem[2648] = 32'b00000010011000000100110111010000;
   assign mem[2649] = 32'b00000001100110011011111000010000;
   assign mem[2650] = 32'b11101000110111101011011010000000;
   assign mem[2651] = 32'b00001010101110111111010001110000;
   assign mem[2652] = 32'b11110001101101110111100111000000;
   assign mem[2653] = 32'b11111001110110010011010111010000;
   assign mem[2654] = 32'b00000101110111110100101010010000;
   assign mem[2655] = 32'b00001011011100111001111001000000;
   assign mem[2656] = 32'b00010001000111111000101110000000;
   assign mem[2657] = 32'b11111111001001101010111000000000;
   assign mem[2658] = 32'b11111011110001001110011101101000;
   assign mem[2659] = 32'b11110010111100001101100100110000;
   assign mem[2660] = 32'b11111101100010110111011010100100;
   assign mem[2661] = 32'b11111101001100000111010000010000;
   assign mem[2662] = 32'b11111110001010111101000101111110;
   assign mem[2663] = 32'b00000000000101101010111001010110;
   assign mem[2664] = 32'b00000011010000111001111111001100;
   assign mem[2665] = 32'b00000100111100100100100001010000;
   assign mem[2666] = 32'b00000010010011111001011000011100;
   assign mem[2667] = 32'b00000001011000110110101110000110;
   assign mem[2668] = 32'b11111111111111101111011000100111;
   assign mem[2669] = 32'b00000010001010011101111010111100;
   assign mem[2670] = 32'b11111111000101110000000101000000;
   assign mem[2671] = 32'b11111011111100001011011000100000;
   assign mem[2672] = 32'b00000010110011000110011111001100;
   assign mem[2673] = 32'b00000001011000110000001110010110;
   assign mem[2674] = 32'b11110110101111101011100001010000;
   assign mem[2675] = 32'b11111000011100001100000111011000;
   assign mem[2676] = 32'b00001001000100100110010100010000;
   assign mem[2677] = 32'b11111010001110010100100001000000;
   assign mem[2678] = 32'b00000101011001010100011101100000;
   assign mem[2679] = 32'b11111100010100100110001011101000;
   assign mem[2680] = 32'b11111101100000011010011001001000;
   assign mem[2681] = 32'b11111111010011101110000010011001;
   assign mem[2682] = 32'b11111011001011010011100000001000;
   assign mem[2683] = 32'b11111111000011100010000101111000;
   assign mem[2684] = 32'b11111001100000000101000101101000;
   assign mem[2685] = 32'b00000100110110000000011111110000;
   assign mem[2686] = 32'b11111001111000100110001000101000;
   assign mem[2687] = 32'b00000110001011111011010011000000;
   assign mem[2688] = 32'b00000100011001110010100000001000;
   assign mem[2689] = 32'b00000010001111100101111100110100;
   assign mem[2690] = 32'b00000010011011000001110001001100;
   assign mem[2691] = 32'b11111011100001001101110011010000;
   assign mem[2692] = 32'b11111101100111101101110011110000;
   assign mem[2693] = 32'b11111100101010110111110001100000;
   assign mem[2694] = 32'b11111110001000010110010001101000;
   assign mem[2695] = 32'b00000001001011110010010111000010;
   assign mem[2696] = 32'b11111111011010111100101000000110;
   assign mem[2697] = 32'b00000000110010011010011101001001;
   assign mem[2698] = 32'b00000001100111001001111110000110;
   assign mem[2699] = 32'b00000000001000110111001110111110;
   assign mem[2700] = 32'b00001000000100101101001011110000;
   assign mem[2701] = 32'b11111011110011000011110001111000;
   assign mem[2702] = 32'b00000010010010010011001000110000;
   assign mem[2703] = 32'b00000010110000100110010001001100;
   assign mem[2704] = 32'b11110110100111001010001111000000;
   assign mem[2705] = 32'b00000100100010000110101001000000;
   assign mem[2706] = 32'b11111100001001100010111110000100;
   assign mem[2707] = 32'b00001011000010001011000110110000;
   assign mem[2708] = 32'b11111111010111000100100001111100;
   assign mem[2709] = 32'b11111100111000111001110010101000;
   assign mem[2710] = 32'b11111100011001110000110011000100;
   assign mem[2711] = 32'b00001010101100001011101111000000;
   assign mem[2712] = 32'b11101010100110110011111110100000;
   assign mem[2713] = 32'b11100000011111101011010011100000;
   assign mem[2714] = 32'b00001010011010001100000100110000;
   assign mem[2715] = 32'b00001001100001111010010000010000;
   assign mem[2716] = 32'b00000011000100110001000000001100;
   assign mem[2717] = 32'b11110101111011110101100111010000;
   assign mem[2718] = 32'b00001001000101101101001100110000;
   assign mem[2719] = 32'b11101000000101111010110100000000;
   assign mem[2720] = 32'b11111110010111111011000110011010;
   assign mem[2721] = 32'b11111101110000010100110100000100;
   assign mem[2722] = 32'b11101110101100100111111110000000;
   assign mem[2723] = 32'b11101111011101011101000111100000;
   assign mem[2724] = 32'b11111011010011010100110001000000;
   assign mem[2725] = 32'b00001010000010000111100110100000;
   assign mem[2726] = 32'b00000000011111111110001010111000;
   assign mem[2727] = 32'b11110010100000001100101100010000;
   assign mem[2728] = 32'b00000110110000111111001100101000;
   assign mem[2729] = 32'b11111001011100001100111000110000;
   assign mem[2730] = 32'b00000010100100001110011011001000;
   assign mem[2731] = 32'b11101111011000100111111010100000;
   assign mem[2732] = 32'b00000111000010110101111111010000;
   assign mem[2733] = 32'b00000110111010101011011011110000;
   assign mem[2734] = 32'b11110000101011111110100001110000;
   assign mem[2735] = 32'b11111000111100111111010000010000;
   assign mem[2736] = 32'b11111111101010101011011011101110;
   assign mem[2737] = 32'b00000000001110011101010000100111;
   assign mem[2738] = 32'b00000000110101000110110110100110;
   assign mem[2739] = 32'b00000011111101011101000110010000;
   assign mem[2740] = 32'b00000101111111101010111010011000;
   assign mem[2741] = 32'b11111110100111010101000101000110;
   assign mem[2742] = 32'b11111111000111110011100110101111;
   assign mem[2743] = 32'b11111111011010111110001101110101;
   assign mem[2744] = 32'b11111111011001000111100110111101;
   assign mem[2745] = 32'b11111010111101000111000111110000;
   assign mem[2746] = 32'b11110111101010100000011011010000;
   assign mem[2747] = 32'b11111111010010011100011010110110;
   assign mem[2748] = 32'b00000011111011101010011101010000;
   assign mem[2749] = 32'b00000010001100111010000110100100;
   assign mem[2750] = 32'b00000001101011110100000111000000;
   assign mem[2751] = 32'b11111110000011011111010111000110;
   assign mem[2752] = 32'b11110011110011100101100010110000;
   assign mem[2753] = 32'b11111110110000000111101011101100;
   assign mem[2754] = 32'b00000001101011000111001110100110;
   assign mem[2755] = 32'b00000100110101110001001100011000;
   assign mem[2756] = 32'b11111101000100001110001000001100;
   assign mem[2757] = 32'b00000010011110111001010010110100;
   assign mem[2758] = 32'b11111110100010000110110101111110;
   assign mem[2759] = 32'b00000100010100000000101010011000;
   assign mem[2760] = 32'b11111011001110111111111100111000;
   assign mem[2761] = 32'b00000010100011110010001111000000;
   assign mem[2762] = 32'b11111000011010101110000100110000;
   assign mem[2763] = 32'b11110101010101010010100111000000;
   assign mem[2764] = 32'b00000011101101111011111101101100;
   assign mem[2765] = 32'b00000000101000101000111111001010;
   assign mem[2766] = 32'b11111101001101000010101000110000;
   assign mem[2767] = 32'b11111110110101101011010110000010;
   assign mem[2768] = 32'b00000100101000111110000101100000;
   assign mem[2769] = 32'b11111001111000100100001110111000;
   assign mem[2770] = 32'b00000001101101010111101111110000;
   assign mem[2771] = 32'b11111100101010000000000011100000;
   assign mem[2772] = 32'b11111100001100111101111101000000;
   assign mem[2773] = 32'b11111110100010001001101101011110;
   assign mem[2774] = 32'b00000101111011110010111011110000;
   assign mem[2775] = 32'b00001000011101000111100101110000;
   assign mem[2776] = 32'b11111100110111111100100110111100;
   assign mem[2777] = 32'b00000010100010101100111100001000;
   assign mem[2778] = 32'b11111111001000110000111111110100;
   assign mem[2779] = 32'b11111111110011010011100010110101;
   assign mem[2780] = 32'b11111110101000111110001111111000;
   assign mem[2781] = 32'b00000110100110111010111000001000;
   assign mem[2782] = 32'b11101110000011011001001101000000;
   assign mem[2783] = 32'b00000010011011111000010001111000;
   assign mem[2784] = 32'b00000101000011111100000101100000;
   assign mem[2785] = 32'b00000010000001010010010000100000;
   assign mem[2786] = 32'b00000110100001011101110000111000;
   assign mem[2787] = 32'b00000101000010001011110100111000;
   assign mem[2788] = 32'b00000010011011001101111100011100;
   assign mem[2789] = 32'b11110101001000101000101100010000;
   assign mem[2790] = 32'b00000011100111111111100111000000;
   assign mem[2791] = 32'b11110111111101100101000111110000;
   assign mem[2792] = 32'b00000011000000001000110101101100;
   assign mem[2793] = 32'b00000001111010001001001011000110;
   assign mem[2794] = 32'b00000010111001010111111101001100;
   assign mem[2795] = 32'b11110000010000001010011111010000;
   assign mem[2796] = 32'b00000001011110011100111000100010;
   assign mem[2797] = 32'b11111101111000110110001011101100;
   assign mem[2798] = 32'b00000000110111011111000100111111;
   assign mem[2799] = 32'b00000000010100011011001111001011;
   assign mem[2800] = 32'b00000100001011110000001001011000;
   assign mem[2801] = 32'b00000110110001110010001011011000;
   assign mem[2802] = 32'b11111101100110101010100000100100;
   assign mem[2803] = 32'b00000000001110010001001011001101;
   assign mem[2804] = 32'b00000001001010011001010001110100;
   assign mem[2805] = 32'b11101110011110110110100110000000;
   assign mem[2806] = 32'b00000101110111110010111010110000;
   assign mem[2807] = 32'b11111010111001000001100000101000;
   assign mem[2808] = 32'b00000100111110100100011000110000;
   assign mem[2809] = 32'b11110110101010110110111101100000;
   assign mem[2810] = 32'b11111010110000000100000101111000;
   assign mem[2811] = 32'b00000110101110001011100110101000;
   assign mem[2812] = 32'b00000100010000101101010101001000;
   assign mem[2813] = 32'b00000011110100100001010100010100;
   assign mem[2814] = 32'b11111100101101000100101100100100;
   assign mem[2815] = 32'b11111101100111011011110101010100;
   assign mem[2816] = 32'b11111110010000001100111000011000;
   assign mem[2817] = 32'b00000001001110101110100101110100;
   assign mem[2818] = 32'b00000110001110001100001010000000;
   assign mem[2819] = 32'b11111101011000100011001110101000;
   assign mem[2820] = 32'b11111111011011000011010110100101;
   assign mem[2821] = 32'b00000011100101110110010000001000;
   assign mem[2822] = 32'b11111100110011111100100110100000;
   assign mem[2823] = 32'b00000011000000001110101111011100;
   assign mem[2824] = 32'b00000000110001011011000000101000;
   assign mem[2825] = 32'b11111001111001101010101000001000;
   assign mem[2826] = 32'b11111111010110010001011011101010;
   assign mem[2827] = 32'b11111100001111001101101100001000;
   assign mem[2828] = 32'b00000000000110011110110011110000;
   assign mem[2829] = 32'b11110111001110010111001001000000;
   assign mem[2830] = 32'b11111101111011010100010010001000;
   assign mem[2831] = 32'b00000111001110001011010010110000;
   assign mem[2832] = 32'b11101000010101100111000001100000;
   assign mem[2833] = 32'b11100010100010010101101001000000;
   assign mem[2834] = 32'b00001110101000101100111101110000;
   assign mem[2835] = 32'b00001011001100101010011111110000;
   assign mem[2836] = 32'b00000101100110001111000000011000;
   assign mem[2837] = 32'b11111111001110000001111010110100;
   assign mem[2838] = 32'b11111100011101100011000111001100;
   assign mem[2839] = 32'b11110010011010001001110101100000;
   assign mem[2840] = 32'b00000100011101111000100010111000;
   assign mem[2841] = 32'b11111110100000110000100111001000;
   assign mem[2842] = 32'b11111010010111100001100010000000;
   assign mem[2843] = 32'b11111110010111101000110101001110;
   assign mem[2844] = 32'b11111011010101101000010110100000;
   assign mem[2845] = 32'b00000101111001101100111000010000;
   assign mem[2846] = 32'b00000000011010010110010000001000;
   assign mem[2847] = 32'b00000100001111101100110010011000;
   assign mem[2848] = 32'b11111100011110001110010110000000;
   assign mem[2849] = 32'b11111011000000010111000110100000;
   assign mem[2850] = 32'b00000011101001011110001111010000;
   assign mem[2851] = 32'b00000001111101110010011101111010;
   assign mem[2852] = 32'b00000000100000100100100001001101;
   assign mem[2853] = 32'b00000000000111011111101010011000;
   assign mem[2854] = 32'b11111101000101000111110111000100;
   assign mem[2855] = 32'b11111111001001000110010110000000;
   assign mem[2856] = 32'b11111111000010110011001110101000;
   assign mem[2857] = 32'b00000010001010111010100100100000;
   assign mem[2858] = 32'b00000000010101001100101111011001;
   assign mem[2859] = 32'b00000001010000000111001100110000;
   assign mem[2860] = 32'b11111000001011100001010000100000;
   assign mem[2861] = 32'b00000101110001101111001100100000;
   assign mem[2862] = 32'b11110111110101100000111011110000;
   assign mem[2863] = 32'b00000110100011001001101000011000;
   assign mem[2864] = 32'b00001001100111110111111001100000;
   assign mem[2865] = 32'b11111010000001100101011111101000;
   assign mem[2866] = 32'b11111111111000000001111110001000;
   assign mem[2867] = 32'b11111011101000101011000010110000;
   assign mem[2868] = 32'b00000101110110000011011000100000;
   assign mem[2869] = 32'b11111001010010010011110010101000;
   assign mem[2870] = 32'b11110111101010111110110001110000;
   assign mem[2871] = 32'b11110100011010100010011001110000;
   assign mem[2872] = 32'b11111100001110111101010001111100;
   assign mem[2873] = 32'b11110011010110010001101111010000;
   assign mem[2874] = 32'b11111100001101010100001011001000;
   assign mem[2875] = 32'b00001000010111100111010000110000;
   assign mem[2876] = 32'b00001101100011010010011110100000;
   assign mem[2877] = 32'b11110001100101101000000110100000;
   assign mem[2878] = 32'b00000000100110110000011111101001;
   assign mem[2879] = 32'b11111001100110001101000110001000;
   assign mem[2880] = 32'b11111100011010001101100010110100;
   assign mem[2881] = 32'b00001001100101111110110001010000;
   assign mem[2882] = 32'b11110111001101001111110010000000;
   assign mem[2883] = 32'b11111011111100100110100101101000;
   assign mem[2884] = 32'b00000101111110000100000001101000;
   assign mem[2885] = 32'b00000001101110000111011010011110;
   assign mem[2886] = 32'b11111100000011101010100110100000;
   assign mem[2887] = 32'b00000100001111111011001101001000;
   assign mem[2888] = 32'b11111010110101010100010001011000;
   assign mem[2889] = 32'b11111011010101101101101110010000;
   assign mem[2890] = 32'b11111000101101001101001001000000;
   assign mem[2891] = 32'b00001010010000101111111110110000;
   assign mem[2892] = 32'b11110000010101011110000011000000;
   assign mem[2893] = 32'b11110000101010000101111000100000;
   assign mem[2894] = 32'b00001101000111011111110010000000;
   assign mem[2895] = 32'b11111110010110110010110100001000;
   assign mem[2896] = 32'b00000001001001101101101010001010;
   assign mem[2897] = 32'b11110111011101000011000000110000;
   assign mem[2898] = 32'b00000110000001000101001011010000;
   assign mem[2899] = 32'b11110110010101000010010110000000;
   assign mem[2900] = 32'b00000010110010010000010010100100;
   assign mem[2901] = 32'b11111001011001110001101000011000;
   assign mem[2902] = 32'b11111010100011011011001010001000;
   assign mem[2903] = 32'b11111100111011110111110001111100;
   assign mem[2904] = 32'b00000011010101001001000100001100;
   assign mem[2905] = 32'b00001000001011111010101000010000;
   assign mem[2906] = 32'b00000010001000100000000111011000;
   assign mem[2907] = 32'b11110100001001111100010111010000;
   assign mem[2908] = 32'b00000001000000001110000101101000;
   assign mem[2909] = 32'b00000001001101100111101001101110;
   assign mem[2910] = 32'b11101001110110101110011100100000;
   assign mem[2911] = 32'b00000101000010101111001011010000;
   assign mem[2912] = 32'b11111001001001100010000100010000;
   assign mem[2913] = 32'b00001000000111101110001110100000;
   assign mem[2914] = 32'b00000000000101001010111110011011;
   assign mem[2915] = 32'b00001000001100001100110101100000;
   assign mem[2916] = 32'b00000101101110110000100101111000;
   assign mem[2917] = 32'b00000001001100101011000001111110;
   assign mem[2918] = 32'b11111111110001011110010110000011;
   assign mem[2919] = 32'b11110100000010001000011011110000;
   assign mem[2920] = 32'b00000110110010001101001101111000;
   assign mem[2921] = 32'b00000011100001101100101111001000;
   assign mem[2922] = 32'b00000010011101111000001010111100;
   assign mem[2923] = 32'b11111111110011010000101110111111;
   assign mem[2924] = 32'b11111101000111111011111011111000;
   assign mem[2925] = 32'b11111101011110011001000100000000;
   assign mem[2926] = 32'b11111111110101101100111010111001;
   assign mem[2927] = 32'b00000001111111000100011100110100;
   assign mem[2928] = 32'b00000011011111111000010100101000;
   assign mem[2929] = 32'b00000001111010111110110000111110;
   assign mem[2930] = 32'b00000010011000111000101000000000;
   assign mem[2931] = 32'b11111110101000010101111010001100;
   assign mem[2932] = 32'b11111111001000110000101111101011;
   assign mem[2933] = 32'b00000100110111010101010001001000;
   assign mem[2934] = 32'b11110111000011110010001000100000;
   assign mem[2935] = 32'b11111100000011001111110101101100;
   assign mem[2936] = 32'b11111101001010000101111110010000;
   assign mem[2937] = 32'b00000000001101111110000000111001;
   assign mem[2938] = 32'b00000011000000101011010011001100;
   assign mem[2939] = 32'b00000001110100111010001001100100;
   assign mem[2940] = 32'b00000101001101010101010011001000;
   assign mem[2941] = 32'b11111101010111001110011010001000;
   assign mem[2942] = 32'b11111101001100110001110001101100;
   assign mem[2943] = 32'b11111100111100100101110100011100;
   assign mem[2944] = 32'b00000000110110011111010011111111;
   assign mem[2945] = 32'b00000101000000010001000000100000;
   assign mem[2946] = 32'b00000001010001000111110111110110;
   assign mem[2947] = 32'b11111011100101110001100010001000;
   assign mem[2948] = 32'b11111100011101111110110101111100;
   assign mem[2949] = 32'b11111101111011000000100100101100;
   assign mem[2950] = 32'b00000001000100011101111111110010;
   assign mem[2951] = 32'b00000110111011001101101000010000;
   assign mem[2952] = 32'b11100110110011110011101001100000;
   assign mem[2953] = 32'b11101011101010101110011100100000;
   assign mem[2954] = 32'b00001100100011100110001000100000;
   assign mem[2955] = 32'b00010010111010000010010001000000;
   assign mem[2956] = 32'b11111110100100001011110011111110;
   assign mem[2957] = 32'b00000011011101010011001111100100;
   assign mem[2958] = 32'b00000000001000011111011011011101;
   assign mem[2959] = 32'b11101111010111010110111010100000;
   assign mem[2960] = 32'b00000101011011101000101010101000;
   assign mem[2961] = 32'b11111010101001111001110101101000;
   assign mem[2962] = 32'b11111011010101110011110110100000;
   assign mem[2963] = 32'b11111011101011011010111111110000;
   assign mem[2964] = 32'b11111001011100111110110001111000;
   assign mem[2965] = 32'b11111010100101110110000101011000;
   assign mem[2966] = 32'b00001000000101001010110111000000;
   assign mem[2967] = 32'b11111000001100010110101101111000;
   assign mem[2968] = 32'b00001100100111011001001001110000;
   assign mem[2969] = 32'b11111100111010010010011010111100;
   assign mem[2970] = 32'b11111100011010100001101101110000;
   assign mem[2971] = 32'b00000000010111001001111010000111;
   assign mem[2972] = 32'b11101000011111000000001100000000;
   assign mem[2973] = 32'b11101111010001000001000110100000;
   assign mem[2974] = 32'b00000001100111110011010011100110;
   assign mem[2975] = 32'b00001001010100011101001101000000;
   assign mem[2976] = 32'b00001100001011011101010101100000;
   assign mem[2977] = 32'b11111010100001110100110001110000;
   assign mem[2978] = 32'b00000011001110100111110011110000;
   assign mem[2979] = 32'b11110011011101000011111001010000;
   assign mem[2980] = 32'b11111100011111011100111000010000;
   assign mem[2981] = 32'b00001001010010101000110100110000;
   assign mem[2982] = 32'b11111000110101100010100010110000;
   assign mem[2983] = 32'b11111001101100101011111100101000;
   assign mem[2984] = 32'b11110010110110100110001011010000;
   assign mem[2985] = 32'b00000110111001001100100001011000;
   assign mem[2986] = 32'b00001000011110010000011110110000;
   assign mem[2987] = 32'b00000011111110001110110010001100;
   assign mem[2988] = 32'b11111010110100101011110011000000;
   assign mem[2989] = 32'b11111011111011101100110011111000;
   assign mem[2990] = 32'b00000000010010011111100100000010;
   assign mem[2991] = 32'b00000010100111011100001001110100;
   assign mem[2992] = 32'b00000101110111011011001111100000;
   assign mem[2993] = 32'b00000101001001100101111110000000;
   assign mem[2994] = 32'b00000000011000110111011110101000;
   assign mem[2995] = 32'b11111010110101010001111110011000;
   assign mem[2996] = 32'b00000000010100100101111100111100;
   assign mem[2997] = 32'b11111011011110101110011001110000;
   assign mem[2998] = 32'b00000001001010110011110110010110;
   assign mem[2999] = 32'b11111001100000111100010010111000;
   assign mem[3000] = 32'b11111111100001010111010010100000;
   assign mem[3001] = 32'b00000001000111010101000001010100;
   assign mem[3002] = 32'b11111001101110111001000000001000;
   assign mem[3003] = 32'b00000010000000110000011111100000;
   assign mem[3004] = 32'b00000100011011001101010101011000;
   assign mem[3005] = 32'b11111110100100001100101000011100;
   assign mem[3006] = 32'b00000101001010010111100110001000;
   assign mem[3007] = 32'b00000010110110111110101001001100;
   assign mem[3008] = 32'b11111110000100010001111000010100;
   assign mem[3009] = 32'b11111111000001111000110101101011;
   assign mem[3010] = 32'b00000110100000010000111001001000;
   assign mem[3011] = 32'b11111001011100101110111111000000;
   assign mem[3012] = 32'b00000111101011010100111010001000;
   assign mem[3013] = 32'b00000100011100110000110001011000;
   assign mem[3014] = 32'b11110100000100001010010100010000;
   assign mem[3015] = 32'b11110110000111110010001101100000;
   assign mem[3016] = 32'b00000010011011100010101011101000;
   assign mem[3017] = 32'b11111011000110011000010010101000;
   assign mem[3018] = 32'b11111111010001111101111011101110;
   assign mem[3019] = 32'b00000011110011100011011110000000;
   assign mem[3020] = 32'b00001010110001011001001000100000;
   assign mem[3021] = 32'b00000001000111100011111011000010;
   assign mem[3022] = 32'b11111011000000111111011010011000;
   assign mem[3023] = 32'b11110010111100110011101010100000;
   assign mem[3024] = 32'b00000111001110101011101011100000;
   assign mem[3025] = 32'b00000101110101010000010111010000;
   assign mem[3026] = 32'b11111100001011000010000110101000;
   assign mem[3027] = 32'b11111110100101000100110110001010;
   assign mem[3028] = 32'b00000101101011011010110101100000;
   assign mem[3029] = 32'b11101110110000100101110001000000;
   assign mem[3030] = 32'b00000000011000100101111111101000;
   assign mem[3031] = 32'b11111011110010100111101101110000;
   assign mem[3032] = 32'b00000001011000110111001010011000;
   assign mem[3033] = 32'b11111011011000100110100100111000;
   assign mem[3034] = 32'b00000010010011010000011001100000;
   assign mem[3035] = 32'b00000010100000010100011000011000;
   assign mem[3036] = 32'b00000001010100100101101000111000;
   assign mem[3037] = 32'b11111100110110011010100101001100;
   assign mem[3038] = 32'b00000010110010100111011000001100;
   assign mem[3039] = 32'b11111101110110101100110001010100;
   assign mem[3040] = 32'b00000011010100001110010010101000;
   assign mem[3041] = 32'b11111011101101001001010001011000;
   assign mem[3042] = 32'b11111000111000011111100010010000;
   assign mem[3043] = 32'b00000011101000111001100011001000;
   assign mem[3044] = 32'b00000101101101010100111110110000;
   assign mem[3045] = 32'b11111111111101100011101000010011;
   assign mem[3046] = 32'b00001000010101000001000100010000;
   assign mem[3047] = 32'b11111010000100101011110011001000;
   assign mem[3048] = 32'b00000000101111111100001001000001;
   assign mem[3049] = 32'b11111011111110010101100110011000;
   assign mem[3050] = 32'b00000001010000111110100111100000;
   assign mem[3051] = 32'b00001000000110000101011000010000;
   assign mem[3052] = 32'b11110100010001111100011100000000;
   assign mem[3053] = 32'b11110011011010001011001000000000;
   assign mem[3054] = 32'b00001000100101010111011001110000;
   assign mem[3055] = 32'b00001001011100100001110110110000;
   assign mem[3056] = 32'b00000000100011010010101011110101;
   assign mem[3057] = 32'b00000010100011010101010111100000;
   assign mem[3058] = 32'b00000001110111001100001101110010;
   assign mem[3059] = 32'b11111001000101000100011001110000;
   assign mem[3060] = 32'b11111011101111101001011011110000;
   assign mem[3061] = 32'b00000100111010110011110001111000;
   assign mem[3062] = 32'b11110110011000110010101001000000;
   assign mem[3063] = 32'b00000010000101000010101010011000;
   assign mem[3064] = 32'b00001110101010100010011011010000;
   assign mem[3065] = 32'b00000101010100100100010111001000;
   assign mem[3066] = 32'b00000100011011001000000011011000;
   assign mem[3067] = 32'b11111011100011111110010010000000;
   assign mem[3068] = 32'b11111101001101010100111001100100;
   assign mem[3069] = 32'b11111010011010101001100100011000;
   assign mem[3070] = 32'b00000000100000101110110100001011;
   assign mem[3071] = 32'b00001001001100100011001111010000;
   assign mem[3072] = 32'b00000010011111000000011111101000;
   assign mem[3073] = 32'b11111000001100100011100110000000;
   assign mem[3074] = 32'b00000110111100101101111011011000;
   assign mem[3075] = 32'b00000110111010000010001011100000;
   assign mem[3076] = 32'b11111111100010111010001111010010;
   assign mem[3077] = 32'b11111100000110111000011011010000;
   assign mem[3078] = 32'b11110101001011001010000101000000;
   assign mem[3079] = 32'b11110100000110110110001101110000;
   assign mem[3080] = 32'b11111110111100010011101111101110;
   assign mem[3081] = 32'b11110100100000001100010000000000;
   assign mem[3082] = 32'b11111110100011110000010011011000;
   assign mem[3083] = 32'b11111011010110110100000110100000;
   assign mem[3084] = 32'b11101100011010001000110010100000;
   assign mem[3085] = 32'b00001000111011101001101010100000;
   assign mem[3086] = 32'b00000100001100110000000001001000;
   assign mem[3087] = 32'b11110110001111001000101010110000;
   assign mem[3088] = 32'b00000101110000000110110110000000;
   assign mem[3089] = 32'b00000011101010101110110111010100;
   assign mem[3090] = 32'b00000000111100101011100011101101;
   assign mem[3091] = 32'b11110111100001000100101000110000;
   assign mem[3092] = 32'b00000001111101010100001100000000;
   assign mem[3093] = 32'b11111111011100100010101001010011;
   assign mem[3094] = 32'b11110111001101111001001110010000;
   assign mem[3095] = 32'b00000100011101011010010100100000;
   assign mem[3096] = 32'b11111111010101110100011011001100;
   assign mem[3097] = 32'b00000101111001001000100010010000;
   assign mem[3098] = 32'b00000010010101011011001011001000;
   assign mem[3099] = 32'b00000001101011111010100110100000;
   assign mem[3100] = 32'b11111000010110011000110100010000;
   assign mem[3101] = 32'b11111101010011101100111101000000;
   assign mem[3102] = 32'b11101011100111000111011111000000;
   assign mem[3103] = 32'b11111110001011011011101011100000;
   assign mem[3104] = 32'b00000101111011101110000101010000;
   assign mem[3105] = 32'b00000101001000001010101010111000;
   assign mem[3106] = 32'b00001101100010001100111101100000;
   assign mem[3107] = 32'b11110101110000101110011110000000;
   assign mem[3108] = 32'b00000001010011010001010101000010;
   assign mem[3109] = 32'b11111010111001011101010101111000;
   assign mem[3110] = 32'b11101101111101000111010100100000;
   assign mem[3111] = 32'b00000101110100010100010110010000;
   assign mem[3112] = 32'b11111011101000010110110101010000;
   assign mem[3113] = 32'b00000101101000010100001111110000;
   assign mem[3114] = 32'b11111111100001011101100110111100;
   assign mem[3115] = 32'b00000100001010011010111001110000;
   assign mem[3116] = 32'b00000010000110100100111110111000;
   assign mem[3117] = 32'b00000100000110101110111000001000;
   assign mem[3118] = 32'b00000000001011111110111100000111;
   assign mem[3119] = 32'b11110110001001100010110111100000;
   assign mem[3120] = 32'b11111000011010110010111001011000;
   assign mem[3121] = 32'b00000110011001010000110110000000;
   assign mem[3122] = 32'b00000011011000111100010011001100;
   assign mem[3123] = 32'b00001000011110110111011110010000;
   assign mem[3124] = 32'b11111111101111100001110101001000;
   assign mem[3125] = 32'b00000000001011111001011100000110;
   assign mem[3126] = 32'b00000000111100010110010000100001;
   assign mem[3127] = 32'b11110110100101110111100101110000;
   assign mem[3128] = 32'b11111111101100000110010101010010;
   assign mem[3129] = 32'b11111101000010010010111001010100;
   assign mem[3130] = 32'b11111111001101101110000101111100;
   assign mem[3131] = 32'b11110100100110011101110110000000;
   assign mem[3132] = 32'b11111110010001010001100000110000;
   assign mem[3133] = 32'b00000010101011111000011001101000;
   assign mem[3134] = 32'b11110000000011001001100110010000;
   assign mem[3135] = 32'b11110101000011000111000001010000;
   assign mem[3136] = 32'b11111110111111001110111001101110;
   assign mem[3137] = 32'b11110110101111010001010111100000;
   assign mem[3138] = 32'b00001010001011011001101111100000;
   assign mem[3139] = 32'b11110000110001010101010111010000;
   assign mem[3140] = 32'b00000001000100011010011001100000;
   assign mem[3141] = 32'b11111101100101011000000011011000;
   assign mem[3142] = 32'b11111011111001110110001101111000;
   assign mem[3143] = 32'b00000000011001100111100111011001;
   assign mem[3144] = 32'b11111111011110000011000011001111;
   assign mem[3145] = 32'b11111101001110001100110001001100;
   assign mem[3146] = 32'b11110111101011001110111101100000;
   assign mem[3147] = 32'b00000001100010010110101010001100;
   assign mem[3148] = 32'b00000011010101001110101011111000;
   assign mem[3149] = 32'b00000000100111000011011000011000;
   assign mem[3150] = 32'b00000110000001100101111111001000;
   assign mem[3151] = 32'b11111100001100001000001011110100;
   assign mem[3152] = 32'b00000001111001011000001000001110;
   assign mem[3153] = 32'b00000001011110111100000100001000;
   assign mem[3154] = 32'b00000010000111110111010011000100;
   assign mem[3155] = 32'b11111101110010011110010011101100;
   assign mem[3156] = 32'b11111011001010011111111010101000;
   assign mem[3157] = 32'b00000100100010001101110100011000;
   assign mem[3158] = 32'b11111101101010010000110101001100;
   assign mem[3159] = 32'b11111011101010000100001100011000;
   assign mem[3160] = 32'b00000001110001001110110000100000;
   assign mem[3161] = 32'b00000110000001101001010110110000;
   assign mem[3162] = 32'b11110100010101100000010010010000;
   assign mem[3163] = 32'b11110110011000001001000110000000;
   assign mem[3164] = 32'b00000111101001100010100101100000;
   assign mem[3165] = 32'b00001100001010000000111010010000;
   assign mem[3166] = 32'b11111110111100110000101010111100;
   assign mem[3167] = 32'b00000001100010011000010110110000;
   assign mem[3168] = 32'b00000001110010101110001100001110;
   assign mem[3169] = 32'b11111000010000110001101101011000;
   assign mem[3170] = 32'b11111010001110110000111100001000;
   assign mem[3171] = 32'b00000011110110110011101011111000;
   assign mem[3172] = 32'b11101101110101101111110010000000;
   assign mem[3173] = 32'b11110010001001001110011110000000;
   assign mem[3174] = 32'b00001000111000000000001110010000;
   assign mem[3175] = 32'b00000110100000100100110010111000;
   assign mem[3176] = 32'b11111010001110010101001101000000;
   assign mem[3177] = 32'b00000100011100001111111110101000;
   assign mem[3178] = 32'b11111110011000110100101000000000;
   assign mem[3179] = 32'b11111111101001010100110110110110;
   assign mem[3180] = 32'b11111001110110000010010110000000;
   assign mem[3181] = 32'b00001100001111011100011101000000;
   assign mem[3182] = 32'b11101001001011101100010001100000;
   assign mem[3183] = 32'b11101001101100001011101101100000;
   assign mem[3184] = 32'b00001011010101100110100000110000;
   assign mem[3185] = 32'b00000000011001000011110101001101;
   assign mem[3186] = 32'b11111001001010010001100011100000;
   assign mem[3187] = 32'b11111100101111100000111111111100;
   assign mem[3188] = 32'b00000110010011011011011010101000;
   assign mem[3189] = 32'b11101010101001111010000101100000;
   assign mem[3190] = 32'b11111110111010110101000101010000;
   assign mem[3191] = 32'b00000101011100110000100111001000;
   assign mem[3192] = 32'b11110111101111000100001111000000;
   assign mem[3193] = 32'b11110101100010001111000101000000;
   assign mem[3194] = 32'b00000010100101101000101100110100;
   assign mem[3195] = 32'b00001011111110110010110000100000;
   assign mem[3196] = 32'b11110111111110010111111010100000;
   assign mem[3197] = 32'b11111111110001110111001011100011;
   assign mem[3198] = 32'b11111110001111110111011000010000;
   assign mem[3199] = 32'b11111001000111100110110111101000;
   assign mem[3200] = 32'b00000001010111000011011101110000;
   assign mem[3201] = 32'b11111000011101111010110100010000;
   assign mem[3202] = 32'b11111010000110110111000111010000;
   assign mem[3203] = 32'b11111111110000110101100101100000;
   assign mem[3204] = 32'b11111110011111000111011101110100;
   assign mem[3205] = 32'b11111111100101110100000001001000;
   assign mem[3206] = 32'b11111110010110110100111110100100;
   assign mem[3207] = 32'b00000000010010111010000010100011;
   assign mem[3208] = 32'b00000101000101101010100000000000;
   assign mem[3209] = 32'b00000101000010000010011110111000;
   assign mem[3210] = 32'b11110110101010000000110110100000;
   assign mem[3211] = 32'b11111001111100111100000100110000;
   assign mem[3212] = 32'b11111110101110010001101000100000;
   assign mem[3213] = 32'b00000011000000001100101111010000;
   assign mem[3214] = 32'b00000100011100010000010100101000;
   assign mem[3215] = 32'b11111100110010101110000010000000;
   assign mem[3216] = 32'b11111111110110101110111101001000;
   assign mem[3217] = 32'b00001100011111011010100111010000;
   assign mem[3218] = 32'b00000011011010101110011000010100;
   assign mem[3219] = 32'b11111101110111000001101001100000;
   assign mem[3220] = 32'b11111100011010001101000101001000;
   assign mem[3221] = 32'b11111100000110010111111100111100;
   assign mem[3222] = 32'b11101111101001111010111001100000;
   assign mem[3223] = 32'b11110101001101110000001001010000;
   assign mem[3224] = 32'b00001101111010101010111010010000;
   assign mem[3225] = 32'b11111101101100100101010010100100;
   assign mem[3226] = 32'b11110111110100101000011100110000;
   assign mem[3227] = 32'b00001011111000011100100111010000;
   assign mem[3228] = 32'b00000110101010011111001011010000;
   assign mem[3229] = 32'b11110100011111000100000111000000;
   assign mem[3230] = 32'b11111100011110001100011101001100;
   assign mem[3231] = 32'b11111011101000011110010011000000;
   assign mem[3232] = 32'b00000010000001001001110011101100;
   assign mem[3233] = 32'b00000101111101001101000110011000;
   assign mem[3234] = 32'b11111110101000100000011001100000;
   assign mem[3235] = 32'b11111000000110110101000000000000;
   assign mem[3236] = 32'b11111010010000001101011101010000;
   assign mem[3237] = 32'b00000000110000111100010110111000;
   assign mem[3238] = 32'b11111111001011000100110000010000;
   assign mem[3239] = 32'b11110101010110001111001011010000;
   assign mem[3240] = 32'b11111101101000011111010111110000;
   assign mem[3241] = 32'b11111101100011111000111110101000;
   assign mem[3242] = 32'b00000101100110010001101000000000;
   assign mem[3243] = 32'b00001010110010110110101000110000;
   assign mem[3244] = 32'b11111010100010110100001100111000;
   assign mem[3245] = 32'b11110100101010100100110000110000;
   assign mem[3246] = 32'b00000100001100000110110101100000;
   assign mem[3247] = 32'b00000011000100110100110110001100;
   assign mem[3248] = 32'b11111001110001101011011011001000;
   assign mem[3249] = 32'b11110011011000101101111011110000;
   assign mem[3250] = 32'b00000000101011111001010001110100;
   assign mem[3251] = 32'b11111111111010010010011000100111;
   assign mem[3252] = 32'b00000101010111110001110110111000;
   assign mem[3253] = 32'b11110011100110001010011000000000;
   assign mem[3254] = 32'b11110111000101101101010010100000;
   assign mem[3255] = 32'b11111010011000011010111000110000;
   assign mem[3256] = 32'b00000101000001101101011101111000;
   assign mem[3257] = 32'b11111111100010010001011101111001;
   assign mem[3258] = 32'b00000000110110011010000010010010;
   assign mem[3259] = 32'b00001010101111100011100000100000;
   assign mem[3260] = 32'b11111011001001010101001011011000;
   assign mem[3261] = 32'b00000001011110100010000110100000;
   assign mem[3262] = 32'b11111110101100110001110001110010;
   assign mem[3263] = 32'b00000000110110010111110011100110;
   assign mem[3264] = 32'b11111000100111111010111101010000;
   assign mem[3265] = 32'b11111110101101111010010010111000;
   assign mem[3266] = 32'b00000110000110000001110011110000;
   assign mem[3267] = 32'b11111000101100100001101100011000;
   assign mem[3268] = 32'b00001000010000000111000001110000;
   assign mem[3269] = 32'b11111111110010111011100011000000;
   assign mem[3270] = 32'b11111010101111011001111111010000;
   assign mem[3271] = 32'b11101111110101010011101010100000;
   assign mem[3272] = 32'b00000111010000000101110110100000;
   assign mem[3273] = 32'b00000010100011101011110010110000;
   assign mem[3274] = 32'b11111101010000001110100000111100;
   assign mem[3275] = 32'b11101000110111011001000111100000;
   assign mem[3276] = 32'b11111110111011001101111010111110;
   assign mem[3277] = 32'b11111011011010100000001000011000;
   assign mem[3278] = 32'b00000000000110111000100001101111;
   assign mem[3279] = 32'b00000011100011010111100010011000;
   assign mem[3280] = 32'b00000110000010010111100101111000;
   assign mem[3281] = 32'b11111101000110001011001110000000;
   assign mem[3282] = 32'b00000011011101001100001011001000;
   assign mem[3283] = 32'b11111010110011100000011010011000;
   assign mem[3284] = 32'b00000001100110100110001000101010;
   assign mem[3285] = 32'b11101111110001101111010110000000;
   assign mem[3286] = 32'b11111110010100011001000010001100;
   assign mem[3287] = 32'b00001101111011001000001101110000;
   assign mem[3288] = 32'b11111111011001111001000011000111;
   assign mem[3289] = 32'b11111010101011110111100000110000;
   assign mem[3290] = 32'b00000001101001001110100100110000;
   assign mem[3291] = 32'b11111010001010000011111110001000;
   assign mem[3292] = 32'b11111011011000011000001011100000;
   assign mem[3293] = 32'b11111010111101100101000110110000;
   assign mem[3294] = 32'b11111110110101101000001100010100;
   assign mem[3295] = 32'b00000010010000000100100110000000;
   assign mem[3296] = 32'b00000100010101011101001110001000;
   assign mem[3297] = 32'b00000001110010111011101000010000;
   assign mem[3298] = 32'b11111111000101001100000010001100;
   assign mem[3299] = 32'b00000001101011000110101000111100;
   assign mem[3300] = 32'b00000100011111101110000001110000;
   assign mem[3301] = 32'b11111011001100000111111101010000;
   assign mem[3302] = 32'b11111100110110010100011101101100;
   assign mem[3303] = 32'b00000000001110000100001000111001;
   assign mem[3304] = 32'b11111010011000010100110110000000;
   assign mem[3305] = 32'b11111111010000101000100100101111;
   assign mem[3306] = 32'b11111101000111111000101000111000;
   assign mem[3307] = 32'b11111111010010110001110000001110;
   assign mem[3308] = 32'b00000001000101001000000100110000;
   assign mem[3309] = 32'b00000000001001001010011011100100;
   assign mem[3310] = 32'b11110110110101011100101101010000;
   assign mem[3311] = 32'b00000101001101110111001011010000;
   assign mem[3312] = 32'b11110110111100001101101001110000;
   assign mem[3313] = 32'b00000000100110010000101101100110;
   assign mem[3314] = 32'b00000110011001110100000001100000;
   assign mem[3315] = 32'b00000110101100011000110001110000;
   assign mem[3316] = 32'b11111000101011100001100100000000;
   assign mem[3317] = 32'b00000111000101110011110111000000;
   assign mem[3318] = 32'b00000011001110110001101100111100;
   assign mem[3319] = 32'b11110111010111011010111111110000;
   assign mem[3320] = 32'b00000101111100100011111100001000;
   assign mem[3321] = 32'b11111111100010010101110010101010;
   assign mem[3322] = 32'b00001011010100011011011110010000;
   assign mem[3323] = 32'b00000101101100111101001101001000;
   assign mem[3324] = 32'b11111111111101100000010000101110;
   assign mem[3325] = 32'b11101001101111010011111000100000;
   assign mem[3326] = 32'b11110110110000011010100000010000;
   assign mem[3327] = 32'b00001010111100011001010011000000;
   assign mem[3328] = 32'b00000011111010111101110101110100;
   assign mem[3329] = 32'b11111000000001010011010010001000;
   assign mem[3330] = 32'b00001001001101100100011111000000;
   assign mem[3331] = 32'b00000000101111100010100011101001;
   assign mem[3332] = 32'b00000110101010101010101011100000;
   assign mem[3333] = 32'b11111110101111101011011001000100;
   assign mem[3334] = 32'b00000010000101111101010111001100;
   assign mem[3335] = 32'b11110111100100100000011101010000;
   assign mem[3336] = 32'b11111011111110010111110001100000;
   assign mem[3337] = 32'b00001010100101101100001001010000;
   assign mem[3338] = 32'b11111011111110010111010111011000;
   assign mem[3339] = 32'b11110101100110111110001011000000;
   assign mem[3340] = 32'b00000000010101011101111111101000;
   assign mem[3341] = 32'b11111010100110111010001100100000;
   assign mem[3342] = 32'b11110100010001110010100110110000;
   assign mem[3343] = 32'b00000000100111101110110010000001;
   assign mem[3344] = 32'b00000100000110101010100011100000;
   assign mem[3345] = 32'b11111111011011110010100111001110;
   assign mem[3346] = 32'b11111111000000011111111100110010;
   assign mem[3347] = 32'b00000111011101010100011010001000;
   assign mem[3348] = 32'b00000110111100110011010101001000;
   assign mem[3349] = 32'b00000010011101111100010100101000;
   assign mem[3350] = 32'b00000100000000100111001001100000;
   assign mem[3351] = 32'b11111100011000011100100110111000;
   assign mem[3352] = 32'b11111100011001001111111101011000;
   assign mem[3353] = 32'b11111011000101010001011010010000;
   assign mem[3354] = 32'b11111110010001100101110101111000;
   assign mem[3355] = 32'b00000001111010000111100100101010;
   assign mem[3356] = 32'b00000010101101110111010110000100;
   assign mem[3357] = 32'b11111111011010101011001111000010;
   assign mem[3358] = 32'b00000001100101010100101010000000;
   assign mem[3359] = 32'b00000001111010110101110110100100;
   assign mem[3360] = 32'b11110001100110011001111001110000;
   assign mem[3361] = 32'b11111101010101010001101001111100;
   assign mem[3362] = 32'b00000010110000110100110000001100;
   assign mem[3363] = 32'b00000101010100000110001000110000;
   assign mem[3364] = 32'b11110011101101110100010000110000;
   assign mem[3365] = 32'b11101011011011001110010001100000;
   assign mem[3366] = 32'b11111110001100010001101110110100;
   assign mem[3367] = 32'b00000010011011111101111001010000;
   assign mem[3368] = 32'b11111110011101101010100000101000;
   assign mem[3369] = 32'b11111000111101101011110100111000;
   assign mem[3370] = 32'b00000100110110011001000111001000;
   assign mem[3371] = 32'b00000000101101101101010001011101;
   assign mem[3372] = 32'b11110110111000011101110000010000;
   assign mem[3373] = 32'b11111001000011110000011110010000;
   assign mem[3374] = 32'b11111110110010000001101111100010;
   assign mem[3375] = 32'b00000110000100000000101101111000;
   assign mem[3376] = 32'b11111011010110001010011100001000;
   assign mem[3377] = 32'b00000101011111111101111101011000;
   assign mem[3378] = 32'b00000000100011011011111011110100;
   assign mem[3379] = 32'b00000100111100111011100101001000;
   assign mem[3380] = 32'b11110101110000100111100100100000;
   assign mem[3381] = 32'b00000001000010110011101011001000;
   assign mem[3382] = 32'b00000110110000001000100010101000;
   assign mem[3383] = 32'b00000110001100010100001100111000;
   assign mem[3384] = 32'b00001000110100011011000011100000;
   assign mem[3385] = 32'b11110001001101000001011010010000;
   assign mem[3386] = 32'b11110100111110111100010011000000;
   assign mem[3387] = 32'b00000110100100011111000110010000;
   assign mem[3388] = 32'b11111010110000011100100000101000;
   assign mem[3389] = 32'b11110100011000100111011111000000;
   assign mem[3390] = 32'b00001001000101000110001111100000;
   assign mem[3391] = 32'b11111111010101111000111110000010;
   assign mem[3392] = 32'b11111011111011110100101001101000;
   assign mem[3393] = 32'b11111010011010110100010111110000;
   assign mem[3394] = 32'b00000011111011100010010010101100;
   assign mem[3395] = 32'b11110010011000000011111010010000;
   assign mem[3396] = 32'b11111100100100011000110010100100;
   assign mem[3397] = 32'b11111001110011100100101101110000;
   assign mem[3398] = 32'b00001001101010110101001110000000;
   assign mem[3399] = 32'b00000111110110010100101100010000;
   assign mem[3400] = 32'b00000001110011010111011110011000;
   assign mem[3401] = 32'b11111011110011001111010010010000;
   assign mem[3402] = 32'b11110101101011000001000001000000;
   assign mem[3403] = 32'b11110111011011100101110100010000;
   assign mem[3404] = 32'b00000010100100001101101011011000;
   assign mem[3405] = 32'b00000001001000001011001111011110;
   assign mem[3406] = 32'b00000001110101111010010100010100;
   assign mem[3407] = 32'b11111110000110111110100100111100;
   assign mem[3408] = 32'b00000001010011000101001101000110;
   assign mem[3409] = 32'b00000000010011111110011010001010;
   assign mem[3410] = 32'b00001000000110100111011000110000;
   assign mem[3411] = 32'b00000001000001000011111111101010;
   assign mem[3412] = 32'b11111111100000010001001001100101;
   assign mem[3413] = 32'b00001000111001000111000101000000;
   assign mem[3414] = 32'b00000101001111000110100011111000;
   assign mem[3415] = 32'b11101001111111100100000011100000;
   assign mem[3416] = 32'b00000000101100000000010001011001;
   assign mem[3417] = 32'b00000001110010110100000000000100;
   assign mem[3418] = 32'b00000100100011111110100000101000;
   assign mem[3419] = 32'b00000011101111010000010100001000;
   assign mem[3420] = 32'b00000100011111001101111101000000;
   assign mem[3421] = 32'b00000011111101110000111011001000;
   assign mem[3422] = 32'b00000010100001100110100101110000;
   assign mem[3423] = 32'b00000001100011011010101100011100;
   assign mem[3424] = 32'b11110101111101100001000011000000;
   assign mem[3425] = 32'b11111101001001101000010100100100;
   assign mem[3426] = 32'b11111110011010000001001110101110;
   assign mem[3427] = 32'b11111101010100110000100110100100;
   assign mem[3428] = 32'b00000100110101110011101011100000;
   assign mem[3429] = 32'b00001000110111100001110111100000;
   assign mem[3430] = 32'b00001011010000100000111010000000;
   assign mem[3431] = 32'b00000001001011101010011011010110;
   assign mem[3432] = 32'b11111011101000111101000001100000;
   assign mem[3433] = 32'b11110001111100001011111101010000;
   assign mem[3434] = 32'b00000100011100001001111010111000;
   assign mem[3435] = 32'b00000001101011111000100110111110;
   assign mem[3436] = 32'b11111011010011101001101111100000;
   assign mem[3437] = 32'b00000000010101110101101100111011;
   assign mem[3438] = 32'b00000011011000011101111010011000;
   assign mem[3439] = 32'b00000011101101010111001100100100;
   assign mem[3440] = 32'b11111011011111101000111100111000;
   assign mem[3441] = 32'b00000100110001111101010000111000;
   assign mem[3442] = 32'b11111000000001000011010010100000;
   assign mem[3443] = 32'b11110111011100000111001111100000;
   assign mem[3444] = 32'b00000001000010000110111101001000;
   assign mem[3445] = 32'b00000010001001011100011000110000;
   assign mem[3446] = 32'b00000010100110111101000110111000;
   assign mem[3447] = 32'b00000100101110111100001110100000;
   assign mem[3448] = 32'b00000101011100011101100010100000;
   assign mem[3449] = 32'b00000010001010001010010011101100;
   assign mem[3450] = 32'b11111010010001110100111111100000;
   assign mem[3451] = 32'b00001010000100000011111001110000;
   assign mem[3452] = 32'b00000010100100111000010110000000;
   assign mem[3453] = 32'b00000011010011000001111111011100;
   assign mem[3454] = 32'b11111000100000101011001111110000;
   assign mem[3455] = 32'b11111101011101010000111010010100;
   assign mem[3456] = 32'b00000110110110110011110001010000;
   assign mem[3457] = 32'b11101011101110011101100110000000;
   assign mem[3458] = 32'b11110111101110100011101111000000;
   assign mem[3459] = 32'b00000010001000101011100110000000;
   assign mem[3460] = 32'b11110001001011010111110011100000;
   assign mem[3461] = 32'b00000110110011001110001111101000;
   assign mem[3462] = 32'b11110010001100011100111100010000;
   assign mem[3463] = 32'b11111010101100000110111101001000;
   assign mem[3464] = 32'b11111110010010001001110100110100;
   assign mem[3465] = 32'b00001100011001011101110111100000;
   assign mem[3466] = 32'b00001101110011110010110010000000;
   assign mem[3467] = 32'b11111110010010111111010100001010;
   assign mem[3468] = 32'b11110101100010010100110111100000;
   assign mem[3469] = 32'b11110001000101011110100111010000;
   assign mem[3470] = 32'b00000011010100111000010100100100;
   assign mem[3471] = 32'b11111001011110010001011000011000;
   assign mem[3472] = 32'b11111111101100011001011000100100;
   assign mem[3473] = 32'b11111100011110001010111111110000;
   assign mem[3474] = 32'b00000001001110011010000101011000;
   assign mem[3475] = 32'b11111101011010110100110010010100;
   assign mem[3476] = 32'b00000001110111001000100110101000;
   assign mem[3477] = 32'b00000000111111101100100101101010;
   assign mem[3478] = 32'b00000000010100101111010001000111;
   assign mem[3479] = 32'b00000011011100000110010110111100;
   assign mem[3480] = 32'b00000000010110001011100111010111;
   assign mem[3481] = 32'b11111010100101110011000010011000;
   assign mem[3482] = 32'b11111110111010110000111000100000;
   assign mem[3483] = 32'b00000000000001001010010010100100;
   assign mem[3484] = 32'b11111100010110001000111110101000;
   assign mem[3485] = 32'b11111001001001001111011001101000;
   assign mem[3486] = 32'b00000010101100001111111000010100;
   assign mem[3487] = 32'b00000001010011101001100001111100;
   assign mem[3488] = 32'b00000000000110010111100010011101;
   assign mem[3489] = 32'b00000100011110111101000010100000;
   assign mem[3490] = 32'b11111111101000100100001000001101;
   assign mem[3491] = 32'b00000100100111011001001110100000;
   assign mem[3492] = 32'b11111111100111000000011111011011;
   assign mem[3493] = 32'b11111110111011110101001101010100;
   assign mem[3494] = 32'b00000011111011101100011100000100;
   assign mem[3495] = 32'b11110110011001000101000001000000;
   assign mem[3496] = 32'b11111101011010111000110000101100;
   assign mem[3497] = 32'b00000111010010101111111101000000;
   assign mem[3498] = 32'b00000011011011111011000110011100;
   assign mem[3499] = 32'b11111011000000100011010111011000;
   assign mem[3500] = 32'b00000000010001101111011100000111;
   assign mem[3501] = 32'b00000001011000110000111110100000;
   assign mem[3502] = 32'b11111010100011110010111011110000;
   assign mem[3503] = 32'b00000000100000011011010101111101;
   assign mem[3504] = 32'b00000010011010000101000110100100;
   assign mem[3505] = 32'b11110001110111001010001101010000;
   assign mem[3506] = 32'b00000101111011011001000101011000;
   assign mem[3507] = 32'b00000100001001000000011000000000;
   assign mem[3508] = 32'b11111011110000100010010100100000;
   assign mem[3509] = 32'b11111101000111110010111110001100;
   assign mem[3510] = 32'b11111000110111001110011100010000;
   assign mem[3511] = 32'b00000110101101000111100111100000;
   assign mem[3512] = 32'b00000110001111011000100001011000;
   assign mem[3513] = 32'b00000101111001001100000001101000;
   assign mem[3514] = 32'b11111111101011110000001110001110;
   assign mem[3515] = 32'b11110111000101101011110111100000;
   assign mem[3516] = 32'b11111110001010001010010101000000;
   assign mem[3517] = 32'b00000110011010111011001011001000;
   assign mem[3518] = 32'b00000010100010101111010100100000;
   assign mem[3519] = 32'b11110100010100011100110100110000;
   assign mem[3520] = 32'b00000111001111000100001010010000;
   assign mem[3521] = 32'b11111010011100011100011111111000;
   assign mem[3522] = 32'b00000001001001100001100110011010;
   assign mem[3523] = 32'b11111101101010111001010011000100;
   assign mem[3524] = 32'b11110101111010001000110101100000;
   assign mem[3525] = 32'b11111010100011000000011000010000;
   assign mem[3526] = 32'b00000001101111111101000001100100;
   assign mem[3527] = 32'b11111110010000101110111000000100;
   assign mem[3528] = 32'b11111110101110100110111011100000;
   assign mem[3529] = 32'b00001000001000100111000110110000;
   assign mem[3530] = 32'b00000010111000111000100100111100;
   assign mem[3531] = 32'b11110110000000100010100010000000;
   assign mem[3532] = 32'b11111001010010111100010011110000;
   assign mem[3533] = 32'b11111001010110000100000011101000;
   assign mem[3534] = 32'b11111101101001110100000001001100;
   assign mem[3535] = 32'b11111110010000011011110101100000;
   assign mem[3536] = 32'b00000001010100000100111100001010;
   assign mem[3537] = 32'b11111001001110100010010110010000;
   assign mem[3538] = 32'b11111111011010001110010011010100;
   assign mem[3539] = 32'b00001000110010001111110010110000;
   assign mem[3540] = 32'b11110101101101001010000111010000;
   assign mem[3541] = 32'b00000100100111011100101011110000;
   assign mem[3542] = 32'b11111011001110101100011111000000;
   assign mem[3543] = 32'b00000010111110011011010000110100;
   assign mem[3544] = 32'b11111100110110101111010001111000;
   assign mem[3545] = 32'b11110110110000101000010000110000;
   assign mem[3546] = 32'b11111100000100111110010011100000;
   assign mem[3547] = 32'b00000100100101001110100001100000;
   assign mem[3548] = 32'b00001010001010001000000111010000;
   assign mem[3549] = 32'b11110101000000110111010001100000;
   assign mem[3550] = 32'b11111101000000101001001010001000;
   assign mem[3551] = 32'b11111100011111000001000101110100;
   assign mem[3552] = 32'b00000101000001101100001000100000;
   assign mem[3553] = 32'b11111011110010001011111101100000;
   assign mem[3554] = 32'b00000001001110011110110001000000;
   assign mem[3555] = 32'b11111000100111011011001011010000;
   assign mem[3556] = 32'b00000010100000110011110000100000;
   assign mem[3557] = 32'b11111010101110010100111110110000;
   assign mem[3558] = 32'b00000101101110100100001110001000;
   assign mem[3559] = 32'b00000000111011000011011001100010;
   assign mem[3560] = 32'b11110010101111000000110011000000;
   assign mem[3561] = 32'b11111111101110000001111000110010;
   assign mem[3562] = 32'b00000101111101100000111100010000;
   assign mem[3563] = 32'b00000010100011010010011111111000;
   assign mem[3564] = 32'b00000000101011101001110000011000;
   assign mem[3565] = 32'b11101100101011001111010000000000;
   assign mem[3566] = 32'b11110111100111011100000101110000;
   assign mem[3567] = 32'b00010001101010111001000111000000;
   assign mem[3568] = 32'b11111101111110000101010101100100;
   assign mem[3569] = 32'b11110010011011101010110111100000;
   assign mem[3570] = 32'b00000011101100111001011101010100;
   assign mem[3571] = 32'b00000101001001101110011111110000;
   assign mem[3572] = 32'b11111011001100111110011011101000;
   assign mem[3573] = 32'b11110110110001110011010100010000;
   assign mem[3574] = 32'b11111111010000100001001100000010;
   assign mem[3575] = 32'b11111110001101000010100010101100;
   assign mem[3576] = 32'b00000011011110110011100101000000;
   assign mem[3577] = 32'b00001010111000111010011001110000;
   assign mem[3578] = 32'b11111101101111100111100110100000;
   assign mem[3579] = 32'b11111110000111101110010001101010;
   assign mem[3580] = 32'b11111110000100001010011111100110;
   assign mem[3581] = 32'b11110100010011111001100000010000;
   assign mem[3582] = 32'b11111110101100010000001010110000;
   assign mem[3583] = 32'b00000011100101000001000111001000;
   assign mem[3584] = 32'b00000101010110010110010011111000;
   assign mem[3585] = 32'b11111110000100110111111100010100;
   assign mem[3586] = 32'b00000010100110011010110011110100;
   assign mem[3587] = 32'b00001010110011111011011111000000;
   assign mem[3588] = 32'b00000111100000101010000011000000;
   assign mem[3589] = 32'b11110000110100010111001000100000;
   assign mem[3590] = 32'b00000100110000101011001101010000;
   assign mem[3591] = 32'b11110100000011111001000100000000;
   assign mem[3592] = 32'b00000010111101100101110110000000;
   assign mem[3593] = 32'b00000001011010100110101100111110;
   assign mem[3594] = 32'b00000111010000000110110011011000;
   assign mem[3595] = 32'b11110010001111101111111011100000;
   assign mem[3596] = 32'b00000000110100000100110010010100;
   assign mem[3597] = 32'b11111100101000010110110111101000;
   assign mem[3598] = 32'b11111101010111101000001011110100;
   assign mem[3599] = 32'b11111100001110100010110000000000;
   assign mem[3600] = 32'b11111011011011011110111101110000;
   assign mem[3601] = 32'b11111111100011101000100010010111;
   assign mem[3602] = 32'b11110011101110110001101011100000;
   assign mem[3603] = 32'b11111111010011111010001011011111;
   assign mem[3604] = 32'b00000111000000011101101011111000;
   assign mem[3605] = 32'b11111101101110111110100110110100;
   assign mem[3606] = 32'b11111010111110001111011011110000;
   assign mem[3607] = 32'b11111110010111000101101001101110;
   assign mem[3608] = 32'b00001011000101010111010010110000;
   assign mem[3609] = 32'b00000010101111100000111110001100;
   assign mem[3610] = 32'b11110010111101100010111111010000;
   assign mem[3611] = 32'b11110111110010001101011000010000;
   assign mem[3612] = 32'b00000110110010001111100001100000;
   assign mem[3613] = 32'b00000010101111100101111000100000;
   assign mem[3614] = 32'b11110100010111111000001010100000;
   assign mem[3615] = 32'b11110000001110000100111111110000;
   assign mem[3616] = 32'b00000001111100100001000110001110;
   assign mem[3617] = 32'b00000000101100010011001011110000;
   assign mem[3618] = 32'b11110110101111001000011001000000;
   assign mem[3619] = 32'b11110001000101100011010010100000;
   assign mem[3620] = 32'b11110110001001010101110110000000;
   assign mem[3621] = 32'b11111110111111110111101111000100;
   assign mem[3622] = 32'b00000001011101101110001000101000;
   assign mem[3623] = 32'b00000101110111010011100101011000;
   assign mem[3624] = 32'b11110011110010000100110010110000;
   assign mem[3625] = 32'b11110111000011101110011010010000;
   assign mem[3626] = 32'b11111110001110101011001010011010;
   assign mem[3627] = 32'b00000101101101100100010111100000;
   assign mem[3628] = 32'b00000001000011110000110100010010;
   assign mem[3629] = 32'b11111011101001011100100001111000;
   assign mem[3630] = 32'b11111000100110010001100001110000;
   assign mem[3631] = 32'b00000011010111010101101011010100;
   assign mem[3632] = 32'b11111011001100110101000001100000;
   assign mem[3633] = 32'b00000011010111000101001001001100;
   assign mem[3634] = 32'b00000100101111001100001011111000;
   assign mem[3635] = 32'b11111010100011100010011111100000;
   assign mem[3636] = 32'b00001100111100000100101011010000;
   assign mem[3637] = 32'b00000000010111010101000100110101;
   assign mem[3638] = 32'b11111110100000110100011111001110;
   assign mem[3639] = 32'b11111001001101000110101001111000;
   assign mem[3640] = 32'b11111111111111011101001011101001;
   assign mem[3641] = 32'b11111111010101011001001111100101;
   assign mem[3642] = 32'b11110100011111000000111100010000;
   assign mem[3643] = 32'b11111111111000110011010000000101;
   assign mem[3644] = 32'b00000010110111111001111000101000;
   assign mem[3645] = 32'b00000000100110111010001100011111;
   assign mem[3646] = 32'b11111010110110100000111011110000;
   assign mem[3647] = 32'b00000011111101010111100001001100;
   assign mem[3648] = 32'b00000110010110011011001001110000;
   assign mem[3649] = 32'b11111100000000110100100101000100;
   assign mem[3650] = 32'b00000011010010011101011011000000;
   assign mem[3651] = 32'b00000000011111100110101000110001;
   assign mem[3652] = 32'b11111011010110110100110110011000;
   assign mem[3653] = 32'b11111111011101011110001110011001;
   assign mem[3654] = 32'b00000110111101000111000000010000;
   assign mem[3655] = 32'b11111011001001001001100010110000;
   assign mem[3656] = 32'b00000000101000000101001101010011;
   assign mem[3657] = 32'b11111110110001111100111110110010;
   assign mem[3658] = 32'b11111110000111101111000110010000;
   assign mem[3659] = 32'b11111101011110101110101000100000;
   assign mem[3660] = 32'b11111111111110101000011101111111;
   assign mem[3661] = 32'b11111011001111000001001100111000;
   assign mem[3662] = 32'b11111100010001111101100010111100;
   assign mem[3663] = 32'b11111101011000010010000000011000;
   assign mem[3664] = 32'b00000000101011010011011111111101;
   assign mem[3665] = 32'b00000010110001111100100100100000;
   assign mem[3666] = 32'b00000010100011011000100000001000;
   assign mem[3667] = 32'b00000000100010101100101101010010;
   assign mem[3668] = 32'b11111101011000100111101011000100;
   assign mem[3669] = 32'b00000010010110001111111000011000;
   assign mem[3670] = 32'b11111111100100100001000010111011;
   assign mem[3671] = 32'b11111100101101100111100111100000;
   assign mem[3672] = 32'b11111011101110000110111101100000;
   assign mem[3673] = 32'b11111111001110101011011101011010;
   assign mem[3674] = 32'b11111100010101101101000110110000;
   assign mem[3675] = 32'b11111111101100011011101000001001;
   assign mem[3676] = 32'b11111101111101110101100101101000;
   assign mem[3677] = 32'b00000000101110111000100011101000;
   assign mem[3678] = 32'b11111100110000110111001100110000;
   assign mem[3679] = 32'b11111111010011101111000100010101;
   assign mem[3680] = 32'b11111001100100100100011100011000;
   assign mem[3681] = 32'b00000000000001110111101000101011;
   assign mem[3682] = 32'b00000000010001101100101111000000;
   assign mem[3683] = 32'b00000000000110110001111011100010;
   assign mem[3684] = 32'b11111011110110111011101110000000;
   assign mem[3685] = 32'b11111010010110001110000101100000;
   assign mem[3686] = 32'b11111110101001001101110001001110;
   assign mem[3687] = 32'b00000101100010001101000000000000;
   assign mem[3688] = 32'b00000001001011010000010001111110;
   assign mem[3689] = 32'b11110111010011110000101010000000;
   assign mem[3690] = 32'b00000111110101000010100101111000;
   assign mem[3691] = 32'b11111111000000000111111000001010;
   assign mem[3692] = 32'b11111000111100111000111001000000;
   assign mem[3693] = 32'b11111101001010000000111001001100;
   assign mem[3694] = 32'b11111100100100110010111000110000;
   assign mem[3695] = 32'b11111111011010010100101011110011;
   assign mem[3696] = 32'b00000010111111010110110110111000;
   assign mem[3697] = 32'b11111111111000010100010001100000;
   assign mem[3698] = 32'b00000000101001000100010000001101;
   assign mem[3699] = 32'b00000010111000001101111000101000;
   assign mem[3700] = 32'b00000100101111001101110011100000;
   assign mem[3701] = 32'b11111101000111100010111011111100;
   assign mem[3702] = 32'b00000010011101110000110010010000;
   assign mem[3703] = 32'b11111111110110011111111110010001;
   assign mem[3704] = 32'b11111000000010101101001101010000;
   assign mem[3705] = 32'b11111010110110110111111110101000;
   assign mem[3706] = 32'b00000010101111011111110111110000;
   assign mem[3707] = 32'b11111100110010111011100111110100;
   assign mem[3708] = 32'b00000011000001011110011111111100;
   assign mem[3709] = 32'b00001001001001010001010101100000;
   assign mem[3710] = 32'b11111110010100110101101010000100;
   assign mem[3711] = 32'b11111110100101110101011011000000;
   assign mem[3712] = 32'b11111111100011000101001110101011;
   assign mem[3713] = 32'b00000001100000001010110110001100;
   assign mem[3714] = 32'b11111111010001001101101100110110;
   assign mem[3715] = 32'b00000000101100011011011110101110;
   assign mem[3716] = 32'b11111110111000110111001000111110;
   assign mem[3717] = 32'b00000010001110100001001011111100;
   assign mem[3718] = 32'b00000010100100100110001110100000;
   assign mem[3719] = 32'b11111011001100101101011100011000;
   assign mem[3720] = 32'b11110100010000110011010011100000;
   assign mem[3721] = 32'b11111000011001001111100100001000;
   assign mem[3722] = 32'b11111111010100110101110100010110;
   assign mem[3723] = 32'b00000011111110010000010101011000;
   assign mem[3724] = 32'b11111001101000110110111100100000;
   assign mem[3725] = 32'b11111100010110100000101010010100;
   assign mem[3726] = 32'b11111001111000011011000001101000;
   assign mem[3727] = 32'b00000111101001101111110011100000;
   assign mem[3728] = 32'b00000001010011001011001010011000;
   assign mem[3729] = 32'b11111101100010101110011111101100;
   assign mem[3730] = 32'b00000000100010111010001101011111;
   assign mem[3731] = 32'b11111000001111000110010101110000;
   assign mem[3732] = 32'b11111100000100001110001101110100;
   assign mem[3733] = 32'b11111110110011100001100011000100;
   assign mem[3734] = 32'b00000011101011110110101011000100;
   assign mem[3735] = 32'b11110001000110011000010011010000;
   assign mem[3736] = 32'b11111110000111100101100010101000;
   assign mem[3737] = 32'b00000110011011010101011001011000;
   assign mem[3738] = 32'b00001011110101000110011101110000;
   assign mem[3739] = 32'b11111111011101101111000001111000;
   assign mem[3740] = 32'b11111000110110110000111001000000;
   assign mem[3741] = 32'b11111100101010101100010110010100;
   assign mem[3742] = 32'b00000011011110010000011001100100;
   assign mem[3743] = 32'b00000011101001000110000110001000;
   assign mem[3744] = 32'b11110010101011110000110101110000;
   assign mem[3745] = 32'b11111011110000000001010010011000;
   assign mem[3746] = 32'b11110110010111001101011101110000;
   assign mem[3747] = 32'b00000010110110111010101001001100;
   assign mem[3748] = 32'b00000011000010100001100000111000;
   assign mem[3749] = 32'b11111110000010011010001100110100;
   assign mem[3750] = 32'b00000001100001101001111001100010;
   assign mem[3751] = 32'b11111111000011100000000101110101;
   assign mem[3752] = 32'b11111101011111000010000101000100;
   assign mem[3753] = 32'b11111111010111001000011100001110;
   assign mem[3754] = 32'b11111010100101111111011100111000;
   assign mem[3755] = 32'b11111100100110010111011011011100;
   assign mem[3756] = 32'b00000110110001000110110110111000;
   assign mem[3757] = 32'b11111111110000100010001111010000;
   assign mem[3758] = 32'b00000011111100110011100010000100;
   assign mem[3759] = 32'b00000100010100000001101110101000;
   assign mem[3760] = 32'b00000001101001010011001110001110;
   assign mem[3761] = 32'b11111111101110010100001101010011;
   assign mem[3762] = 32'b11111101011010011111001110001100;
   assign mem[3763] = 32'b00000000111011001100100000001001;
   assign mem[3764] = 32'b00000011000101101011010010011000;
   assign mem[3765] = 32'b11111011110000100110111010101000;
   assign mem[3766] = 32'b00000011110101110011010010001000;
   assign mem[3767] = 32'b11111101011100101110101010000100;
   assign mem[3768] = 32'b00000010011111000101000100111100;
   assign mem[3769] = 32'b11111100101011111010100011101100;
   assign mem[3770] = 32'b11111100101100100111010111111000;
   assign mem[3771] = 32'b00000100010010110110111001111000;
   assign mem[3772] = 32'b11111011100110100101111110000000;
   assign mem[3773] = 32'b00000000110001010110100100101101;
   assign mem[3774] = 32'b00001000010100000010111010110000;
   assign mem[3775] = 32'b11111010000101111111110011010000;
   assign mem[3776] = 32'b11111000000001100011101110000000;
   assign mem[3777] = 32'b11111111001001110010101010000011;
   assign mem[3778] = 32'b00000100100010010010110000110000;
   assign mem[3779] = 32'b11111010111000010000000100101000;
   assign mem[3780] = 32'b00000011110001111011101111000000;
   assign mem[3781] = 32'b11111101111110010111101011010100;
   assign mem[3782] = 32'b00000011111010011011100010011100;
   assign mem[3783] = 32'b11111010101101101010010010000000;
   assign mem[3784] = 32'b00000011110001100111110000100100;
   assign mem[3785] = 32'b11110011110101101000001101000000;
   assign mem[3786] = 32'b11111111011000111011111001001100;
   assign mem[3787] = 32'b00000101011111100100011011111000;
   assign mem[3788] = 32'b11111100001110000111001100000100;
   assign mem[3789] = 32'b11111100001110001111000110111100;
   assign mem[3790] = 32'b00000001011110111111011110111110;
   assign mem[3791] = 32'b11111011011100110001010111000000;
   assign mem[3792] = 32'b11111011100001000110101011010000;
   assign mem[3793] = 32'b11111101110110011101110101100000;
   assign mem[3794] = 32'b00000110000100100101000101001000;
   assign mem[3795] = 32'b11111001101110010110111101010000;
   assign mem[3796] = 32'b11111111101000110000100000001100;
   assign mem[3797] = 32'b00000110100011110010100111010000;
   assign mem[3798] = 32'b11111111111110111001010011000100;
   assign mem[3799] = 32'b11111111101000100010010010001111;
   assign mem[3800] = 32'b00000011101000011111000100110100;
   assign mem[3801] = 32'b00000000011110011101101111000001;
   assign mem[3802] = 32'b11111111000000110011010110100000;
   assign mem[3803] = 32'b11111101001001101100010001010100;
   assign mem[3804] = 32'b00000010010100101101111001101100;
   assign mem[3805] = 32'b11110111100111010010010100100000;
   assign mem[3806] = 32'b11111111100111101001010100011011;
   assign mem[3807] = 32'b00000001010101011110010110110010;
   assign mem[3808] = 32'b11111111011110101010110001111010;
   assign mem[3809] = 32'b00000001010011110111011110011100;
   assign mem[3810] = 32'b00000001101101101010111100111000;
   assign mem[3811] = 32'b11111111110000111111001000011100;
   assign mem[3812] = 32'b11111001010110110101101011110000;
   assign mem[3813] = 32'b11111101100000110101100110010100;
   assign mem[3814] = 32'b11111100001000011101010000100000;
   assign mem[3815] = 32'b00000011001111011010011111101100;
   assign mem[3816] = 32'b00000011001011111001110001101000;
   assign mem[3817] = 32'b11111100010110101100100011111100;
   assign mem[3818] = 32'b00000011100110111111000011001000;
   assign mem[3819] = 32'b00000011000110100101010110101000;
   assign mem[3820] = 32'b00000010011100101000011110111100;
   assign mem[3821] = 32'b11111010111001110110001111110000;
   assign mem[3822] = 32'b11111010101011100101100000000000;
   assign mem[3823] = 32'b11111011000010111010001110000000;
   assign mem[3824] = 32'b00000011101001011111111110111100;
   assign mem[3825] = 32'b11111111101010011001001110001111;
   assign mem[3826] = 32'b00000110101111011110011010000000;
   assign mem[3827] = 32'b00000001000100110010011001111000;
   assign mem[3828] = 32'b00000011001011101010110111101000;
   assign mem[3829] = 32'b00000000000010111111010010110100;
   assign mem[3830] = 32'b00000000100000011000000000010001;
   assign mem[3831] = 32'b11110111010001010001111010000000;
   assign mem[3832] = 32'b11111010110111011101000000001000;
   assign mem[3833] = 32'b11111000100011111000110001011000;
   assign mem[3834] = 32'b00000010111100010111111110111100;
   assign mem[3835] = 32'b00000001100110010001101101101010;
   assign mem[3836] = 32'b00000100011111110110100000010000;
   assign mem[3837] = 32'b00000010110110001110101110001000;
   assign mem[3838] = 32'b11111101001010101110101001111100;
   assign mem[3839] = 32'b00000011100011000000011001111000;
   assign mem[3840] = 32'b11110101001001001011111100110000;
   assign mem[3841] = 32'b11111110000011110101100101000000;
   assign mem[3842] = 32'b00000000111010000101101010000010;
   assign mem[3843] = 32'b11111111011101110010011111010100;
   assign mem[3844] = 32'b11111001110000000100011110101000;
   assign mem[3845] = 32'b11111110011101000101001000001000;
   assign mem[3846] = 32'b11110001011000000110101010100000;
   assign mem[3847] = 32'b11111100101000101000000010110000;
   assign mem[3848] = 32'b00001011101010011010010111000000;
   assign mem[3849] = 32'b00001011100000101011101001000000;
   assign mem[3850] = 32'b11110110001101110001110111000000;
   assign mem[3851] = 32'b00000100010010110001111100110000;
   assign mem[3852] = 32'b11111100101011110011001011010100;
   assign mem[3853] = 32'b00000001110110100110010101000010;
   assign mem[3854] = 32'b00001100011000100110100100110000;
   assign mem[3855] = 32'b11111111001011100011001000100001;
   assign mem[3856] = 32'b11111010110001000000110110100000;
   assign mem[3857] = 32'b00001101001110111000110110100000;
   assign mem[3858] = 32'b11111011101010010101010000110000;
   assign mem[3859] = 32'b11100100011110100010111010100000;
   assign mem[3860] = 32'b11110010010101101111011100010000;
   assign mem[3861] = 32'b00000011110111000100011100000000;
   assign mem[3862] = 32'b11111110001000010110011010010010;
   assign mem[3863] = 32'b11110100101111110011110001010000;
   assign mem[3864] = 32'b00000100010001100110110110111000;
   assign mem[3865] = 32'b11111111101000010111110111010011;
   assign mem[3866] = 32'b11110101010000100000010011000000;
   assign mem[3867] = 32'b00000100101010111100101111110000;
   assign mem[3868] = 32'b00001001101000111000000010000000;
   assign mem[3869] = 32'b00001011110011011101000101010000;
   assign mem[3870] = 32'b11111001111100001010011010000000;
   assign mem[3871] = 32'b00000101100000001101110111100000;
   assign mem[3872] = 32'b00000100000001000001011101011000;
   assign mem[3873] = 32'b00000110110110110101100011011000;
   assign mem[3874] = 32'b11110101000100111100110000010000;
   assign mem[3875] = 32'b11111010100000110101110101111000;
   assign mem[3876] = 32'b11110000011110010111001100110000;
   assign mem[3877] = 32'b00000101100011100000101010000000;
   assign mem[3878] = 32'b11111001000110011011000001101000;
   assign mem[3879] = 32'b11110110111111010011100011000000;
   assign mem[3880] = 32'b11111001000110001101001100011000;
   assign mem[3881] = 32'b00000010100110001001010111110000;
   assign mem[3882] = 32'b00000100100110011011100100110000;
   assign mem[3883] = 32'b00001000010101001001110001100000;
   assign mem[3884] = 32'b11101011101000011111100010000000;
   assign mem[3885] = 32'b11110100111101011010011110100000;
   assign mem[3886] = 32'b00000000010000010110010100111001;
   assign mem[3887] = 32'b00000111100110101101001010000000;
   assign mem[3888] = 32'b11101101000011010011010111000000;
   assign mem[3889] = 32'b11111100000010011000111001000000;
   assign mem[3890] = 32'b11111110010000111111010000110010;
   assign mem[3891] = 32'b11110000010010100111111111100000;
   assign mem[3892] = 32'b00000100000000000010011111001000;
   assign mem[3893] = 32'b11110100010100100111110011000000;
   assign mem[3894] = 32'b00000000001111110011000100010111;
   assign mem[3895] = 32'b00000011000100100111000000100100;
   assign mem[3896] = 32'b00000110001100000110010001010000;
   assign mem[3897] = 32'b11111011101100001001110111011000;
   assign mem[3898] = 32'b00000000101000000101110101001101;
   assign mem[3899] = 32'b00000010100110110000101011011100;
   assign mem[3900] = 32'b11111011001010011011111001001000;
   assign mem[3901] = 32'b11111011110001001111010011101000;
   assign mem[3902] = 32'b11111100000001110110100101010100;
   assign mem[3903] = 32'b11101110011010000111011000100000;
   assign mem[3904] = 32'b00001000101111001110101001110000;
   assign mem[3905] = 32'b00000100010001101110110000000000;
   assign mem[3906] = 32'b00010000100100101000001010000000;
   assign mem[3907] = 32'b11101111000110010000110111100000;
   assign mem[3908] = 32'b11111011111100110111101111011000;
   assign mem[3909] = 32'b00000101000111010101010111110000;
   assign mem[3910] = 32'b11111110000010100100010101101110;
   assign mem[3911] = 32'b11111100001011101001011010101100;
   assign mem[3912] = 32'b00000010110100010000010001111000;
   assign mem[3913] = 32'b00001000101100110010011111110000;
   assign mem[3914] = 32'b11111110010101100101011111110000;
   assign mem[3915] = 32'b11111001100010100011101100001000;
   assign mem[3916] = 32'b00000000010110100010001001000010;
   assign mem[3917] = 32'b11111111001110000100001001001100;
   assign mem[3918] = 32'b00000001000111000111000001010110;
   assign mem[3919] = 32'b00000010000100010000000100001000;
   assign mem[3920] = 32'b11111111011000001100010100111100;
   assign mem[3921] = 32'b00000001011101100000101001111000;
   assign mem[3922] = 32'b00000100001100110011000001011000;
   assign mem[3923] = 32'b00000000100101011110011001101111;
   assign mem[3924] = 32'b11111100101100010100011001011100;
   assign mem[3925] = 32'b11111001110010010000010010001000;
   assign mem[3926] = 32'b11111011111000101110011110111000;
   assign mem[3927] = 32'b00001000100100100111110000110000;
   assign mem[3928] = 32'b11111101011000001111000010101100;
   assign mem[3929] = 32'b11110101101100100010111111010000;
   assign mem[3930] = 32'b11111111011110101010001010001101;
   assign mem[3931] = 32'b11111110111010000110010011010010;
   assign mem[3932] = 32'b11111111001001111100101100101010;
   assign mem[3933] = 32'b11110011000001001110011011100000;
   assign mem[3934] = 32'b00000000000111110101111011101010;
   assign mem[3935] = 32'b00000001111100101101000110111000;
   assign mem[3936] = 32'b00000011101011100101000101000100;
   assign mem[3937] = 32'b00000001000110011000111001000010;
   assign mem[3938] = 32'b00000011000010010000001000111000;
   assign mem[3939] = 32'b00000011010001101110001110110000;
   assign mem[3940] = 32'b00000001101101110111001111111010;
   assign mem[3941] = 32'b00000010100010111111001000100100;
   assign mem[3942] = 32'b11111110100100001011111001100000;
   assign mem[3943] = 32'b11111111101010101010010010110010;
   assign mem[3944] = 32'b11111101100100110100000011110100;
   assign mem[3945] = 32'b11111010100011010110100011101000;
   assign mem[3946] = 32'b11111101110111010100111111000000;
   assign mem[3947] = 32'b00000100101110001001010010100000;
   assign mem[3948] = 32'b00000010110111101010000111100000;
   assign mem[3949] = 32'b00000010100000110100111111100000;
   assign mem[3950] = 32'b11110010010110110100010111010000;
   assign mem[3951] = 32'b00000101011101010111001001100000;
   assign mem[3952] = 32'b11111110000110111101111101111110;
   assign mem[3953] = 32'b11111011010000100111000001110000;
   assign mem[3954] = 32'b11111010101111111010010010111000;
   assign mem[3955] = 32'b11111100101101100100101011111100;
   assign mem[3956] = 32'b11110001111110011110111110110000;
   assign mem[3957] = 32'b00000001111100011101001010100100;
   assign mem[3958] = 32'b00000100100110010001101011101000;
   assign mem[3959] = 32'b00000110001010011010001000001000;
   assign mem[3960] = 32'b11111111101110100110010111010100;
   assign mem[3961] = 32'b11111010001010101010000101001000;
   assign mem[3962] = 32'b00000010101101100011001110111000;
   assign mem[3963] = 32'b11110100010101100101011110000000;
   assign mem[3964] = 32'b00000101101110101011110111011000;
   assign mem[3965] = 32'b11111100111011101101101100100100;
   assign mem[3966] = 32'b11111001010010011011001001101000;
   assign mem[3967] = 32'b00000101000010000110100011011000;
   assign mem[3968] = 32'b00000101101011100001001001110000;
   assign mem[3969] = 32'b00000000100110101010110111001100;
   assign mem[3970] = 32'b00000110000000100100001011101000;
   assign mem[3971] = 32'b00000110101100010111111011110000;
   assign mem[3972] = 32'b00000110111100101110000011111000;
   assign mem[3973] = 32'b11110101010101101011101110100000;
   assign mem[3974] = 32'b11111101000110000011101100010000;
   assign mem[3975] = 32'b11111001101010011110111000111000;
   assign mem[3976] = 32'b11110111001100101101110110000000;
   assign mem[3977] = 32'b00001111010010010001000110100000;
   assign mem[3978] = 32'b11111110101111100000101100011100;
   assign mem[3979] = 32'b11110101101010010001111110100000;
   assign mem[3980] = 32'b11111011110101011011100001000000;
   assign mem[3981] = 32'b11111100011011100000101111011000;
   assign mem[3982] = 32'b11110111110010000010011010000000;
   assign mem[3983] = 32'b11110111111100101010101111110000;
   assign mem[3984] = 32'b00000110101000010110101000010000;
   assign mem[3985] = 32'b00000010011111100001000001010000;
   assign mem[3986] = 32'b11111110011011101101011011001000;
   assign mem[3987] = 32'b11111110100101110101111000101010;
   assign mem[3988] = 32'b00000111100011100110100001111000;
   assign mem[3989] = 32'b00001001101101101011111010110000;
   assign mem[3990] = 32'b11111110001100000000000011111100;
   assign mem[3991] = 32'b11111000111110110011010110111000;
   assign mem[3992] = 32'b11111010011110100101100111001000;
   assign mem[3993] = 32'b11111010100100100011000010111000;
   assign mem[3994] = 32'b00000000011110000001011010110001;
   assign mem[3995] = 32'b00000100001000110111100001111000;
   assign mem[3996] = 32'b00000010100111011111101100011100;
   assign mem[3997] = 32'b00000011101011111110110000001100;
   assign mem[3998] = 32'b00000000100101011010000011001000;
   assign mem[3999] = 32'b00000101000100101011111000101000;
   assign mem[4000] = 32'b11111110110100010001010001000100;
   assign mem[4001] = 32'b00000100100100110100111000100000;
   assign mem[4002] = 32'b11111111010100100001110000010110;
   assign mem[4003] = 32'b00000100111011111100010100100000;
   assign mem[4004] = 32'b11111010110001010001100100001000;
   assign mem[4005] = 32'b11111100101001001000001111010100;
   assign mem[4006] = 32'b11111001110000111111100111101000;
   assign mem[4007] = 32'b00000111011100110101001110000000;
   assign mem[4008] = 32'b11110110010011110101011010000000;
   assign mem[4009] = 32'b11111001110000001100111100000000;
   assign mem[4010] = 32'b00000010111111001011011101001000;
   assign mem[4011] = 32'b00000100110110011001000000110000;
   assign mem[4012] = 32'b00000011101010011010001100001000;
   assign mem[4013] = 32'b11110000100011110111011111100000;
   assign mem[4014] = 32'b11111100010100101101111000110000;
   assign mem[4015] = 32'b00000011110100101010110111110100;
   assign mem[4016] = 32'b11111101100101110101011101100100;
   assign mem[4017] = 32'b11111111100110000101101001011010;
   assign mem[4018] = 32'b11111111101111110101110011101000;
   assign mem[4019] = 32'b00000000011001111110101101101011;
   assign mem[4020] = 32'b11111100110001010110100010110100;
   assign mem[4021] = 32'b11110001111110001100100010010000;
   assign mem[4022] = 32'b00000111001111011000101110001000;
   assign mem[4023] = 32'b11110101010100001000101100000000;
   assign mem[4024] = 32'b11111111010111101000101011011001;
   assign mem[4025] = 32'b00000000101110001110110101101010;
   assign mem[4026] = 32'b11111101100100000011001100110100;
   assign mem[4027] = 32'b00000101111000101111011000001000;
   assign mem[4028] = 32'b11111100010111100000101110010000;
   assign mem[4029] = 32'b00001000000111010001101001000000;
   assign mem[4030] = 32'b00000000001111010101101100011000;
   assign mem[4031] = 32'b11111110110001100100010001010100;
   assign mem[4032] = 32'b11111111001010111100111011000110;
   assign mem[4033] = 32'b11111100101110100100001111001100;
   assign mem[4034] = 32'b00000001000101001011100101110000;
   assign mem[4035] = 32'b11110110101001001111010101000000;
   assign mem[4036] = 32'b00000100011110100010001001101000;
   assign mem[4037] = 32'b11111010101111000110100100001000;
   assign mem[4038] = 32'b11111011110100110000100111100000;
   assign mem[4039] = 32'b00000110101110100011111101011000;
   assign mem[4040] = 32'b00000001000100000100101011000110;
   assign mem[4041] = 32'b11111101000000101010011000001000;
   assign mem[4042] = 32'b11111111100000001011111010101100;
   assign mem[4043] = 32'b11110011000111101111110011100000;
   assign mem[4044] = 32'b00000001111000111001110010000100;
   assign mem[4045] = 32'b00000001110111101010001010101010;
   assign mem[4046] = 32'b00000100100110010110100110111000;
   assign mem[4047] = 32'b00000011001100010000011111101100;
   assign mem[4048] = 32'b00000000111001001101111101100011;
   assign mem[4049] = 32'b00000001101110111110010111001000;
   assign mem[4050] = 32'b11111111100011001110101011000010;
   assign mem[4051] = 32'b11111111111110110010100101111101;
   assign mem[4052] = 32'b11111010010001000010111101001000;
   assign mem[4053] = 32'b00000011100011110011011111101000;
   assign mem[4054] = 32'b11111110101001001101011011011100;
   assign mem[4055] = 32'b11111110110001011000001011001100;
   assign mem[4056] = 32'b11111101110011100000101101011000;
   assign mem[4057] = 32'b00000011101001011010010011100100;
   assign mem[4058] = 32'b11111101011111101010110111010100;
   assign mem[4059] = 32'b00000010110010010111010111010000;
   assign mem[4060] = 32'b11111110001001001010100100101100;
   assign mem[4061] = 32'b11111000111101001010110000100000;
   assign mem[4062] = 32'b11111111011100011101110100111100;
   assign mem[4063] = 32'b00000011111000101110001010001000;
   assign mem[4064] = 32'b00000010101100011101001100001000;
   assign mem[4065] = 32'b11111100011100011111011010101100;
   assign mem[4066] = 32'b00000101000011011110001000110000;
   assign mem[4067] = 32'b11111101101000100101001101110100;
   assign mem[4068] = 32'b00000100110110100101110000001000;
   assign mem[4069] = 32'b00000001010101100010100100001000;
   assign mem[4070] = 32'b00000001011111111011111110110010;
   assign mem[4071] = 32'b00000001000011100110111101001000;
   assign mem[4072] = 32'b11111101111110111100001110100000;
   assign mem[4073] = 32'b11101111011010101001011111000000;
   assign mem[4074] = 32'b00000110110111000101001100111000;
   assign mem[4075] = 32'b00000000010000000100101010010100;
   assign mem[4076] = 32'b11111110000010010001011110011000;
   assign mem[4077] = 32'b00000001110001001000011110101000;
   assign mem[4078] = 32'b00000011100101000110100000001000;
   assign mem[4079] = 32'b00000101101011101000111101101000;
   assign mem[4080] = 32'b11111001111000011010111100110000;
   assign mem[4081] = 32'b00000010010100100100100001000100;
   assign mem[4082] = 32'b11110101001101001001000001100000;
   assign mem[4083] = 32'b11110000011101111011001101010000;
   assign mem[4084] = 32'b00000111110100010011000110011000;
   assign mem[4085] = 32'b00000010000100110111010110110000;
   assign mem[4086] = 32'b11111110011000111110110001101110;
   assign mem[4087] = 32'b00000100111010001101100000100000;
   assign mem[4088] = 32'b00000001010100011110010011001010;
   assign mem[4089] = 32'b00000100010000001011100101111000;
   assign mem[4090] = 32'b11111101101001001110010011111100;
   assign mem[4091] = 32'b11111110011110101011111100001010;
   assign mem[4092] = 32'b11111111010010001101100110111000;
   assign mem[4093] = 32'b11111000011100010110110111111000;
   assign mem[4094] = 32'b00000110010010100111001110100000;
   assign mem[4095] = 32'b11111010000011111000010001110000;
   assign mem[4096] = 32'b00001111010010010111101011100000;
   assign mem[4097] = 32'b11110100100101101010001001100000;
   assign mem[4098] = 32'b11111101010011101110001111010000;
   assign mem[4099] = 32'b11111111000100011010001111101110;
   assign mem[4100] = 32'b11111110101100100110100000111010;
   assign mem[4101] = 32'b11111000101000100110100100010000;
   assign mem[4102] = 32'b11110100110101100011101010000000;
   assign mem[4103] = 32'b11100110110110011101101101100000;
   assign mem[4104] = 32'b00001011100000010010111110110000;
   assign mem[4105] = 32'b00000000111000000100010111010110;
   assign mem[4106] = 32'b00001100010100101100011111010000;
   assign mem[4107] = 32'b11111001100100011101110110110000;
   assign mem[4108] = 32'b11111111000101011011110100001001;
   assign mem[4109] = 32'b00000010011110011100001110000100;
   assign mem[4110] = 32'b00000010100111110001110100101100;
   assign mem[4111] = 32'b11111011000011000011111010010000;
   assign mem[4112] = 32'b11111110001001101110101110110000;
   assign mem[4113] = 32'b11111110100000000010111010000010;
   assign mem[4114] = 32'b00000001101001101001000001100110;
   assign mem[4115] = 32'b00000001001101100110110000010110;
   assign mem[4116] = 32'b00000011110010100110100110000100;
   assign mem[4117] = 32'b11111100110000101100111110111100;
   assign mem[4118] = 32'b00000010011011111100010100111000;
   assign mem[4119] = 32'b00000010001000111000011011010100;
   assign mem[4120] = 32'b11111101100010100101011011101100;
   assign mem[4121] = 32'b00000000011011101001110101011100;
   assign mem[4122] = 32'b11110111010100111110011000010000;
   assign mem[4123] = 32'b11111100110101010101100011001000;
   assign mem[4124] = 32'b00000010111011100011011110101100;
   assign mem[4125] = 32'b11111101011001111100100101101000;
   assign mem[4126] = 32'b00001001011000010111101010100000;
   assign mem[4127] = 32'b00000010110000110000100011000100;
   assign mem[4128] = 32'b00000101011110101101100100000000;
   assign mem[4129] = 32'b00000111100010001111101110001000;
   assign mem[4130] = 32'b00000101000111000000110011101000;
   assign mem[4131] = 32'b11111111111101011100010111010101;
   assign mem[4132] = 32'b00000011010010000101001110111100;
   assign mem[4133] = 32'b00000000001110011011001100101001;
   assign mem[4134] = 32'b11110101100101000111011111010000;
   assign mem[4135] = 32'b11111100010111110101110001101000;
   assign mem[4136] = 32'b11110110000101101010111100000000;
   assign mem[4137] = 32'b00000111110010101001010010000000;
   assign mem[4138] = 32'b11111100001111101001001111000000;
   assign mem[4139] = 32'b11111110001100101110100110110110;
   assign mem[4140] = 32'b00000100111010111110010001000000;
   assign mem[4141] = 32'b11101000100110111000010000100000;
   assign mem[4142] = 32'b00000000100010110000101011001100;
   assign mem[4143] = 32'b11111000100001101011100111101000;
   assign mem[4144] = 32'b00000110111001111110101011111000;
   assign mem[4145] = 32'b00000010011010101011111010001100;
   assign mem[4146] = 32'b00000011111100111001001111001100;
   assign mem[4147] = 32'b00000101110101111110100011010000;
   assign mem[4148] = 32'b11111100100000110010101000011100;
   assign mem[4149] = 32'b11111110010000000010000111001010;
   assign mem[4150] = 32'b11111111111000000100000011101111;
   assign mem[4151] = 32'b00000011011101100010011001111000;
   assign mem[4152] = 32'b00000011111001010110010010010100;
   assign mem[4153] = 32'b00000101001001001000001101111000;
   assign mem[4154] = 32'b11110011001011010101111111110000;
   assign mem[4155] = 32'b00000001001001011101001100101110;
   assign mem[4156] = 32'b11110101101010001100110101100000;
   assign mem[4157] = 32'b00000101011010101111010111000000;
   assign mem[4158] = 32'b11111011011000101010100000000000;
   assign mem[4159] = 32'b00000100001110001010000101000000;
   assign mem[4160] = 32'b00000000001010111000011011001111;
   assign mem[4161] = 32'b11110011100001010011101100110000;
   assign mem[4162] = 32'b00000010110011101100111101000100;
   assign mem[4163] = 32'b11111100101100010110101010010100;
   assign mem[4164] = 32'b11111110011000011001001000110110;
   assign mem[4165] = 32'b11111100011000100111011011011000;
   assign mem[4166] = 32'b11111101011001101100100011100000;
   assign mem[4167] = 32'b11111100101101001010001000101100;
   assign mem[4168] = 32'b00000001000110110010001100011100;
   assign mem[4169] = 32'b00000100101110100011111100101000;
   assign mem[4170] = 32'b00000010000010101001000101000000;
   assign mem[4171] = 32'b11111000100100001001010111000000;
   assign mem[4172] = 32'b00000000010111100100100101100111;
   assign mem[4173] = 32'b11111011011010010010100011111000;
   assign mem[4174] = 32'b00000001000110111010101100110110;
   assign mem[4175] = 32'b11111100101001100010011010011100;
   assign mem[4176] = 32'b00000101001010100011000001101000;
   assign mem[4177] = 32'b00000000111000011111110100101111;
   assign mem[4178] = 32'b00000011001100110000101101001000;
   assign mem[4179] = 32'b00000011001110011110000011101000;
   assign mem[4180] = 32'b00000011100000010111100001100100;
   assign mem[4181] = 32'b00000000011001101100110010000010;
   assign mem[4182] = 32'b11111111000100101001010100000010;
   assign mem[4183] = 32'b11111101101110010111101110110100;
   assign mem[4184] = 32'b11110110001010011111001010010000;
   assign mem[4185] = 32'b11111100000011000000100100010100;
   assign mem[4186] = 32'b11111011110011110011001100011000;
   assign mem[4187] = 32'b00000111101001101010111110001000;
   assign mem[4188] = 32'b00000000010110111111111111011001;
   assign mem[4189] = 32'b00001001111110100011101001000000;
   assign mem[4190] = 32'b00000000111111000101011110110100;
   assign mem[4191] = 32'b11111010001011100100010110101000;
   assign mem[4192] = 32'b11111111110110011100100111101111;
   assign mem[4193] = 32'b11111111001010011001011000111011;
   assign mem[4194] = 32'b00000011000010011001000011110100;
   assign mem[4195] = 32'b00000001000010001101010111100100;
   assign mem[4196] = 32'b00000101111000111100110101110000;
   assign mem[4197] = 32'b11111000000110000101010111000000;
   assign mem[4198] = 32'b11111100110101010001101101011100;
   assign mem[4199] = 32'b00000100111000100011111000011000;
   assign mem[4200] = 32'b11110011111101100010100000100000;
   assign mem[4201] = 32'b11111000001110100011100111110000;
   assign mem[4202] = 32'b00000111000111000110111001011000;
   assign mem[4203] = 32'b11111100101100101100000000110100;
   assign mem[4204] = 32'b00000000101010101011000110101101;
   assign mem[4205] = 32'b11111011101001000111101111010000;
   assign mem[4206] = 32'b11110101011010011001010111000000;
   assign mem[4207] = 32'b00001101000010110011001100010000;
   assign mem[4208] = 32'b00000110010001000110110101001000;
   assign mem[4209] = 32'b11111001011100101010110010011000;
   assign mem[4210] = 32'b00000101011111001010011101001000;
   assign mem[4211] = 32'b11111100111010010000010011111000;
   assign mem[4212] = 32'b11111000011011000101011001100000;
   assign mem[4213] = 32'b00000000001100100001001001010010;
   assign mem[4214] = 32'b00000010110111000001011010000000;
   assign mem[4215] = 32'b00000000101101110100111010001110;
   assign mem[4216] = 32'b11111011111101110111001100011000;
   assign mem[4217] = 32'b00001001000010010110000101100000;
   assign mem[4218] = 32'b00000110001000010000001001011000;
   assign mem[4219] = 32'b11110011110110001110100100110000;
   assign mem[4220] = 32'b00000001010011101101110001100100;
   assign mem[4221] = 32'b11111101011101010010111100111000;
   assign mem[4222] = 32'b11110111011000100111100101000000;
   assign mem[4223] = 32'b11111101010111001110100101001000;
   assign mem[4224] = 32'b00000011100010010011100110111100;
   assign mem[4225] = 32'b00000010111001100100010001110100;
   assign mem[4226] = 32'b11111011111010100100100110101000;
   assign mem[4227] = 32'b00000101011000011110001011000000;
   assign mem[4228] = 32'b00000001111111000000000001000010;
   assign mem[4229] = 32'b11111010011010111010011000001000;
   assign mem[4230] = 32'b11111111011110110001001000000110;
   assign mem[4231] = 32'b11111100100011100101110011101100;
   assign mem[4232] = 32'b00000011111101111110110101010100;
   assign mem[4233] = 32'b00001000000001101111001100110000;
   assign mem[4234] = 32'b11111011111011100011101001101000;
   assign mem[4235] = 32'b11111100111100100100000110011000;
   assign mem[4236] = 32'b00000000000101011010110110000010;
   assign mem[4237] = 32'b00000011001110110111000100111000;
   assign mem[4238] = 32'b11111010011000101010101110111000;
   assign mem[4239] = 32'b11111001001001100111000000010000;
   assign mem[4240] = 32'b11111001100011011100111111000000;
   assign mem[4241] = 32'b00000100001111001100111010100000;
   assign mem[4242] = 32'b00000010100111000001111111001100;
   assign mem[4243] = 32'b11110111100110000100111001110000;
   assign mem[4244] = 32'b11111001110001101110100001100000;
   assign mem[4245] = 32'b00000010100101110011110100111100;
   assign mem[4246] = 32'b11110111000110000010001100010000;
   assign mem[4247] = 32'b11111101001101000111110101000000;
   assign mem[4248] = 32'b00000000110000010100101101101100;
   assign mem[4249] = 32'b00001110100111110000110100100000;
   assign mem[4250] = 32'b00000110011110011001100101010000;
   assign mem[4251] = 32'b11111011000101100000100111110000;
   assign mem[4252] = 32'b00000110001001011111110000111000;
   assign mem[4253] = 32'b00000010011111111001111101011000;
   assign mem[4254] = 32'b11110011100100001010010111000000;
   assign mem[4255] = 32'b11111011100110000111000110111000;
   assign mem[4256] = 32'b11111111010010010011100010001111;
   assign mem[4257] = 32'b00000101111110101000101000010000;
   assign mem[4258] = 32'b11110110110110101110101010000000;
   assign mem[4259] = 32'b11111011111011010101011011010000;
   assign mem[4260] = 32'b11111010001011010110111100010000;
   assign mem[4261] = 32'b00000100101010010111011110100000;
   assign mem[4262] = 32'b00000011110011110100101110011100;
   assign mem[4263] = 32'b00001000100101100101001111010000;
   assign mem[4264] = 32'b11101001110010001111011001000000;
   assign mem[4265] = 32'b11111011000010100110000100110000;
   assign mem[4266] = 32'b11110110100101111010001110100000;
   assign mem[4267] = 32'b00000101111100111010011101100000;
   assign mem[4268] = 32'b00000000001101001110011110111101;
   assign mem[4269] = 32'b00000000010010000101001010001111;
   assign mem[4270] = 32'b11111110011011100000010000011000;
   assign mem[4271] = 32'b11111011111100010101000010111000;
   assign mem[4272] = 32'b11101010100011110010011001000000;
   assign mem[4273] = 32'b11110100101110110101111001000000;
   assign mem[4274] = 32'b00010001011001010011001110000000;
   assign mem[4275] = 32'b11111110011111110100100100100100;
   assign mem[4276] = 32'b00000010001111101101110011101100;
   assign mem[4277] = 32'b00001011111110100011100100100000;
   assign mem[4278] = 32'b11110111011000010100100011110000;
   assign mem[4279] = 32'b11110110111101100101101111010000;
   assign mem[4280] = 32'b11111111101011011001101101111000;
   assign mem[4281] = 32'b11111100000000100100110001100100;
   assign mem[4282] = 32'b11111101000100100100110011101000;
   assign mem[4283] = 32'b11110011000011000101100011010000;
   assign mem[4284] = 32'b00000011100001011011011001111100;
   assign mem[4285] = 32'b00000001110101110000100110011110;
   assign mem[4286] = 32'b00000000011000011001011010010111;
   assign mem[4287] = 32'b11111100011000110010000100100000;
   assign mem[4288] = 32'b00000011110000000001100011100100;
   assign mem[4289] = 32'b00001010000000010101000101100000;
   assign mem[4290] = 32'b00000010011001010101010000100100;
   assign mem[4291] = 32'b11111011111001011011010001000000;
   assign mem[4292] = 32'b11111101001101111001000000011000;
   assign mem[4293] = 32'b11111100010010011000111001011100;
   assign mem[4294] = 32'b00001000100110001000001101100000;
   assign mem[4295] = 32'b11110110110111100101010110110000;
   assign mem[4296] = 32'b11111100011101101100111000100000;
   assign mem[4297] = 32'b00001110011011100111100011010000;
   assign mem[4298] = 32'b00000100101000110011011000100000;
   assign mem[4299] = 32'b11111000000100011011100100111000;
   assign mem[4300] = 32'b11111100001100001001011100000100;
   assign mem[4301] = 32'b11111100010010101010011101000000;
   assign mem[4302] = 32'b00000000011101000110110111101001;
   assign mem[4303] = 32'b11111100111101100001100110000000;
   assign mem[4304] = 32'b11111110010010011010000011101010;
   assign mem[4305] = 32'b00000011001011110110001000101000;
   assign mem[4306] = 32'b00000001110011010010111001110110;
   assign mem[4307] = 32'b11111111111000100001111101001101;
   assign mem[4308] = 32'b00000001010100111011001000101110;
   assign mem[4309] = 32'b00000000010011001001010010001010;
   assign mem[4310] = 32'b11111111010111100110010101000111;
   assign mem[4311] = 32'b00000011011010100110101100000000;
   assign mem[4312] = 32'b11111110011011000111010000000110;
   assign mem[4313] = 32'b00000011010001100001111101101000;
   assign mem[4314] = 32'b11111101010001011000101111011100;
   assign mem[4315] = 32'b11111100001111011101110010101100;
   assign mem[4316] = 32'b11111100111001110101000000110100;
   assign mem[4317] = 32'b00000000100101111010101110010101;
   assign mem[4318] = 32'b11111110111010110010110001000000;
   assign mem[4319] = 32'b11111100110010101011101011100000;
   assign mem[4320] = 32'b00001100011111111100100010100000;
   assign mem[4321] = 32'b11110111010011000110001001100000;
   assign mem[4322] = 32'b00000001100110110111010111100100;
   assign mem[4323] = 32'b00000000000100111101010111001001;
   assign mem[4324] = 32'b11110111001100100110110111010000;
   assign mem[4325] = 32'b00000010110110011010101000000100;
   assign mem[4326] = 32'b00000010011110010001000000010100;
   assign mem[4327] = 32'b00000010111011011111000101000100;
   assign mem[4328] = 32'b00000011011110111100100000111000;
   assign mem[4329] = 32'b11111110000000110001011010100100;
   assign mem[4330] = 32'b00000001111101000000010100001100;
   assign mem[4331] = 32'b11111100000001001001011000000100;
   assign mem[4332] = 32'b11111100011011101100100110110000;
   assign mem[4333] = 32'b11111011001110101001011100001000;
   assign mem[4334] = 32'b00000100001000111100100110011000;
   assign mem[4335] = 32'b11111111100100010110100100100100;
   assign mem[4336] = 32'b00000010111011011100111110110000;
   assign mem[4337] = 32'b00000001100010010011100101000010;
   assign mem[4338] = 32'b00000001000001001111000111100000;
   assign mem[4339] = 32'b00000010101100001100111011000100;
   assign mem[4340] = 32'b00000000110100000010110001011111;
   assign mem[4341] = 32'b11111111110010000110100111001010;
   assign mem[4342] = 32'b11111001111100011010110100101000;
   assign mem[4343] = 32'b00000001000111010100100110011000;
   assign mem[4344] = 32'b00000011011100111010010101000000;
   assign mem[4345] = 32'b11111010001100010111010111010000;
   assign mem[4346] = 32'b00000001101101110001110010111100;
   assign mem[4347] = 32'b11111110000010100100000111001010;
   assign mem[4348] = 32'b00000010000011010111010100101100;
   assign mem[4349] = 32'b00000101010000100010100101000000;
   assign mem[4350] = 32'b11111010000011001001011000010000;
   assign mem[4351] = 32'b00000000101101010100000000010011;
   assign mem[4352] = 32'b00000010001010100011111111001100;
   assign mem[4353] = 32'b11111111110010011001011100110101;
   assign mem[4354] = 32'b11111111101100010100110110011100;
   assign mem[4355] = 32'b00000000110100110001101011011111;
   assign mem[4356] = 32'b11110100111011000001111001110000;
   assign mem[4357] = 32'b00000001110000000100111100111100;
   assign mem[4358] = 32'b00000010000111110000110001011100;
   assign mem[4359] = 32'b11111111001000111111001111111010;
   assign mem[4360] = 32'b00000010111101011001101101010000;
   assign mem[4361] = 32'b00000001000000111100001110000110;
   assign mem[4362] = 32'b00000011001001010001000110011000;
   assign mem[4363] = 32'b00000100100000010001110001110000;
   assign mem[4364] = 32'b11110111111011001110101100100000;
   assign mem[4365] = 32'b11111101000010010010011001111000;
   assign mem[4366] = 32'b11110100111010111100011101110000;
   assign mem[4367] = 32'b00000010000000101011111100000000;
   assign mem[4368] = 32'b11111100001010101111001101111100;
   assign mem[4369] = 32'b00000001110000001111101010010000;
   assign mem[4370] = 32'b00000000010011010111010010100100;
   assign mem[4371] = 32'b11110110101100110111111010010000;
   assign mem[4372] = 32'b00000011001110000001000011111100;
   assign mem[4373] = 32'b11111101111010100001000001011100;
   assign mem[4374] = 32'b11110111001011010100001111110000;
   assign mem[4375] = 32'b00000000110101010101110100010010;
   assign mem[4376] = 32'b11111000100000001001110100011000;
   assign mem[4377] = 32'b00000101001001110100000011111000;
   assign mem[4378] = 32'b00000010001110001000100011001000;
   assign mem[4379] = 32'b00001000100010101011110000000000;
   assign mem[4380] = 32'b11111110011110001000010001111110;
   assign mem[4381] = 32'b11111011110010111001000110000000;
   assign mem[4382] = 32'b00000010010001101101110010000100;
   assign mem[4383] = 32'b00000010101111100000000011010100;
   assign mem[4384] = 32'b11111010101100011101101111100000;
   assign mem[4385] = 32'b11111100001011110100100001101100;
   assign mem[4386] = 32'b11110110111100111011010011000000;
   assign mem[4387] = 32'b00000010100100010000011101000000;
   assign mem[4388] = 32'b11111010101011100101011011110000;
   assign mem[4389] = 32'b00000010000011111100111110011100;
   assign mem[4390] = 32'b00000001011011001011110100101010;
   assign mem[4391] = 32'b11110011010011110011001011110000;
   assign mem[4392] = 32'b11111101111100101111100011001000;
   assign mem[4393] = 32'b11111101001001001100111100101000;
   assign mem[4394] = 32'b00000011100110110001010101001000;
   assign mem[4395] = 32'b00000000110001000111010000011100;
   assign mem[4396] = 32'b00001000101011100100010000100000;
   assign mem[4397] = 32'b11110111111000101011111110110000;
   assign mem[4398] = 32'b11111011000001001101000001100000;
   assign mem[4399] = 32'b00000111101000110011111000101000;
   assign mem[4400] = 32'b00000000110111010101001001011000;
   assign mem[4401] = 32'b11111110100000111100011100111100;
   assign mem[4402] = 32'b11111101111000010001110101010100;
   assign mem[4403] = 32'b00000101011010011001110000011000;
   assign mem[4404] = 32'b00001010010111010000000101100000;
   assign mem[4405] = 32'b11111110011100110000100111110110;
   assign mem[4406] = 32'b00000000011010100001010110000010;
   assign mem[4407] = 32'b00000100101101001111100101001000;
   assign mem[4408] = 32'b11111110100100101001111001111000;
   assign mem[4409] = 32'b11101111110101011100110110000000;
   assign mem[4410] = 32'b11110110110001001101110111010000;
   assign mem[4411] = 32'b00000010110010010111111000111000;
   assign mem[4412] = 32'b11111111001100100010011110011100;
   assign mem[4413] = 32'b00000011100110110101111101011000;
   assign mem[4414] = 32'b11111101111110010001000110101100;
   assign mem[4415] = 32'b00000110011101010000100100100000;
   assign mem[4416] = 32'b11101111110011110010010001000000;
   assign mem[4417] = 32'b00000100000000001001010001101000;
   assign mem[4418] = 32'b00000010100111000111000110110000;
   assign mem[4419] = 32'b11111000001011100111110011110000;
   assign mem[4420] = 32'b00000011100000000110010101011100;
   assign mem[4421] = 32'b00000010010101010100010101001000;
   assign mem[4422] = 32'b11111101010000000110011000111000;
   assign mem[4423] = 32'b11111101100111011110010010000000;
   assign mem[4424] = 32'b00000010111001001111110011101000;
   assign mem[4425] = 32'b11111110010100010001010011111010;
   assign mem[4426] = 32'b11111110110011011001001100010110;
   assign mem[4427] = 32'b00001111001010100110101000010000;
   assign mem[4428] = 32'b11111011000110011101001000011000;
   assign mem[4429] = 32'b11110010111011010110110011000000;
   assign mem[4430] = 32'b00000001111100100111100000000110;
   assign mem[4431] = 32'b11111011111001001001110101100000;
   assign mem[4432] = 32'b11111101000110000011001011101000;
   assign mem[4433] = 32'b11111000001101001100111000100000;
   assign mem[4434] = 32'b00001001000100001111001010100000;
   assign mem[4435] = 32'b00000001000000000111011101110100;
   assign mem[4436] = 32'b00000010100000000101110010010000;
   assign mem[4437] = 32'b00000101111110110011000101100000;
   assign mem[4438] = 32'b11110110110001110000011101100000;
   assign mem[4439] = 32'b11111010001111100011000011001000;
   assign mem[4440] = 32'b11111101010000100100000110010000;
   assign mem[4441] = 32'b11111010110101010110101010111000;
   assign mem[4442] = 32'b11111110100100100101011101011000;
   assign mem[4443] = 32'b00000011110000011001101001001000;
   assign mem[4444] = 32'b11111111101110000001110010000010;
   assign mem[4445] = 32'b11111101011010010000110000010100;
   assign mem[4446] = 32'b11111101000001000101001000000100;
   assign mem[4447] = 32'b11111011101010000011010001110000;
   assign mem[4448] = 32'b11111101010011010011110101100000;
   assign mem[4449] = 32'b00000001100111100110001111011000;
   assign mem[4450] = 32'b00000011110000100010000001111100;
   assign mem[4451] = 32'b11111000111011111000000100110000;
   assign mem[4452] = 32'b11111011101001110000100111011000;
   assign mem[4453] = 32'b11110111100110010100001101000000;
   assign mem[4454] = 32'b00000000101010111110110000010010;
   assign mem[4455] = 32'b00000000101001010000001101011010;
   assign mem[4456] = 32'b00000000111000000101010110100011;
   assign mem[4457] = 32'b11111101010100111111000111100000;
   assign mem[4458] = 32'b00000010011000011011010001100100;
   assign mem[4459] = 32'b00000100111111010110100010010000;
   assign mem[4460] = 32'b00000001000001110011001101011000;
   assign mem[4461] = 32'b00000000001110100001011100010010;
   assign mem[4462] = 32'b00000000010010100000101100010100;
   assign mem[4463] = 32'b11110110011101101001101011100000;
   assign mem[4464] = 32'b00000110001101111001110001101000;
   assign mem[4465] = 32'b00000110001110111001001111111000;
   assign mem[4466] = 32'b00000010000100110011000111100000;
   assign mem[4467] = 32'b00000011010110011000100010001100;
   assign mem[4468] = 32'b00000011000001000000110111010100;
   assign mem[4469] = 32'b11111110101100010001001011011010;
   assign mem[4470] = 32'b00000100110100010010011001001000;
   assign mem[4471] = 32'b11111010011010111001110110011000;
   assign mem[4472] = 32'b11111100110100110101000101000100;
   assign mem[4473] = 32'b11110010100100111000011100110000;
   assign mem[4474] = 32'b00000011010110111111011100111000;
   assign mem[4475] = 32'b00000100010110110001110001011000;
   assign mem[4476] = 32'b00000011001100010111001100001100;
   assign mem[4477] = 32'b00001001010011010111000001000000;
   assign mem[4478] = 32'b00000001011100001110101111001110;
   assign mem[4479] = 32'b00000011101111110001011101111100;
   assign mem[4480] = 32'b11111010001110101101111101011000;
   assign mem[4481] = 32'b11101101111111001101000010000000;
   assign mem[4482] = 32'b11111111101010000110111001000101;
   assign mem[4483] = 32'b11111101101010011001010001111000;
   assign mem[4484] = 32'b00000011001110010111010011100100;
   assign mem[4485] = 32'b11111110001100000101101111111000;
   assign mem[4486] = 32'b00000100100111011110101011000000;
   assign mem[4487] = 32'b11111101010001111001110001010000;
   assign mem[4488] = 32'b00000011101100110111001111110000;
   assign mem[4489] = 32'b00000100011010001111001010110000;
   assign mem[4490] = 32'b11111101000010010110111110000100;
   assign mem[4491] = 32'b00001100011011111000000111000000;
   assign mem[4492] = 32'b00000111010100101001010011001000;
   assign mem[4493] = 32'b11111000001001111110010110011000;
   assign mem[4494] = 32'b00000110010111011010111011010000;
   assign mem[4495] = 32'b11111110110110011001000100111110;
   assign mem[4496] = 32'b11111001000110001010100100111000;
   assign mem[4497] = 32'b00000000001101011010000011011011;
   assign mem[4498] = 32'b11101011111101011000111100100000;
   assign mem[4499] = 32'b11100011100101010101110010100000;
   assign mem[4500] = 32'b00000101110011000111101000111000;
   assign mem[4501] = 32'b00000000110101010111111010000010;
   assign mem[4502] = 32'b00000001000001111010101100100010;
   assign mem[4503] = 32'b11111101011111111100000001010000;
   assign mem[4504] = 32'b11110011000110000000110110100000;
   assign mem[4505] = 32'b11111100110011101111001000101000;
   assign mem[4506] = 32'b11111111011110011110101011110011;
   assign mem[4507] = 32'b11111011011010011010101010110000;
   assign mem[4508] = 32'b00001001000011000010001111000000;
   assign mem[4509] = 32'b00000101111010010100101110101000;
   assign mem[4510] = 32'b11111001000111011101111010110000;
   assign mem[4511] = 32'b00000011111010010110010100101000;
   assign mem[4512] = 32'b00000100010001111010100000110000;
   assign mem[4513] = 32'b00000111000100010100101111101000;
   assign mem[4514] = 32'b11111100000111000000100011100100;
   assign mem[4515] = 32'b11111101101101011010101011100100;
   assign mem[4516] = 32'b11110110000110010000011101100000;
   assign mem[4517] = 32'b00001001010001100010000110000000;
   assign mem[4518] = 32'b11111011100011001011101001111000;
   assign mem[4519] = 32'b11111110100100101101110000001110;
   assign mem[4520] = 32'b11111100010100101101011111011100;
   assign mem[4521] = 32'b00000000111010001000100001010101;
   assign mem[4522] = 32'b00000111100111111101000010000000;
   assign mem[4523] = 32'b11111111101100001110110011111001;
   assign mem[4524] = 32'b11110100011011111110000001010000;
   assign mem[4525] = 32'b11111100101000111010011101101000;
   assign mem[4526] = 32'b11111100101111001000100100100100;
   assign mem[4527] = 32'b00000111111011110110001100000000;
   assign mem[4528] = 32'b11110011101110101100000111110000;
   assign mem[4529] = 32'b00000000011011010111101000011101;
   assign mem[4530] = 32'b00000010111110000011010000111100;
   assign mem[4531] = 32'b11111011000110101011110111001000;
   assign mem[4532] = 32'b11111010111101111000001110100000;
   assign mem[4533] = 32'b11111011010110101111111001110000;
   assign mem[4534] = 32'b00000011010100011100110011010100;
   assign mem[4535] = 32'b11111100110000110110110000111100;
   assign mem[4536] = 32'b00000001110100011000111100000110;
   assign mem[4537] = 32'b11111010001010001100011100101000;
   assign mem[4538] = 32'b00000100010101000110101110001000;
   assign mem[4539] = 32'b00000101011011100011111010010000;
   assign mem[4540] = 32'b00000001011100101101111100001000;
   assign mem[4541] = 32'b11111110101000010011011001001110;
   assign mem[4542] = 32'b11111100000100011100001000001100;
   assign mem[4543] = 32'b11111001011011101001100000110000;
   assign mem[4544] = 32'b00000111011010111010111110110000;
   assign mem[4545] = 32'b00000011011001000001000100100100;
   assign mem[4546] = 32'b00001001001010101101010110010000;
   assign mem[4547] = 32'b11111110110111011111000110000100;
   assign mem[4548] = 32'b11111101011110000010000100000100;
   assign mem[4549] = 32'b11110110110110111001010101100000;
   assign mem[4550] = 32'b00000011000001000111111101100100;
   assign mem[4551] = 32'b11111111010111010001001110000011;
   assign mem[4552] = 32'b00001000100101110111001100000000;
   assign mem[4553] = 32'b11111100010101100011000101010000;
   assign mem[4554] = 32'b00000010100111110000010011110100;
   assign mem[4555] = 32'b11111010111110010100001000001000;
   assign mem[4556] = 32'b00000101001000011010111100010000;
   assign mem[4557] = 32'b11111111010100000000011001101100;
   assign mem[4558] = 32'b00000000000111110010110101100011;
   assign mem[4559] = 32'b00000010111010001010010101100100;
   assign mem[4560] = 32'b00000110110001111101100110000000;
   assign mem[4561] = 32'b11111000011101010110011010000000;
   assign mem[4562] = 32'b00001000010001010100101101110000;
   assign mem[4563] = 32'b11111111110110001000001110111011;
   assign mem[4564] = 32'b11111000000001000100111001001000;
   assign mem[4565] = 32'b11111001000010001111100010011000;
   assign mem[4566] = 32'b11111000100101101000110011010000;
   assign mem[4567] = 32'b00000110000111000100110111110000;
   assign mem[4568] = 32'b11111110111010110010011000001110;
   assign mem[4569] = 32'b11111110101110011110010110100010;
   assign mem[4570] = 32'b11110111111111011100100100100000;
   assign mem[4571] = 32'b00000011010110101011000101000100;
   assign mem[4572] = 32'b00000011010001111011000000010000;
   assign mem[4573] = 32'b11110011110011010100101111000000;
   assign mem[4574] = 32'b11111101111111000001100000100100;
   assign mem[4575] = 32'b00000110100010011101111110011000;
   assign mem[4576] = 32'b00000010110000101011001101000000;
   assign mem[4577] = 32'b11111111111000001001111111010101;
   assign mem[4578] = 32'b11111111010011111010000000001110;
   assign mem[4579] = 32'b00000010110111110100111111010000;
   assign mem[4580] = 32'b11111100000100001111001001011100;
   assign mem[4581] = 32'b00000001100010010100001000011000;
   assign mem[4582] = 32'b11111101011100100011000011101000;
   assign mem[4583] = 32'b00000001111100110001001101010110;
   assign mem[4584] = 32'b11111111101011000100010110101100;
   assign mem[4585] = 32'b11111011010111111100101001001000;
   assign mem[4586] = 32'b11111010111011001110111100010000;
   assign mem[4587] = 32'b00000010101001111000001101001100;
   assign mem[4588] = 32'b11111111111011000011000111001100;
   assign mem[4589] = 32'b00000000101111101001001100100100;
   assign mem[4590] = 32'b00000100110000100001000010101000;
   assign mem[4591] = 32'b11111101000101000001111101101100;
   assign mem[4592] = 32'b00000010011101000001100001110100;
   assign mem[4593] = 32'b11111100111000100111100010100100;
   assign mem[4594] = 32'b11110011000100100001100111100000;
   assign mem[4595] = 32'b00000011010000001110110000111000;
   assign mem[4596] = 32'b11110000100010010011110010010000;
   assign mem[4597] = 32'b00000100111011111100001111101000;
   assign mem[4598] = 32'b00001001001100101001010001010000;
   assign mem[4599] = 32'b00001000101110001001010110100000;
   assign mem[4600] = 32'b11111000101001010100000011101000;
   assign mem[4601] = 32'b11110000100110000111001101000000;
   assign mem[4602] = 32'b00000010001111110001010010101100;
   assign mem[4603] = 32'b11111111010010101010100111010111;
   assign mem[4604] = 32'b00000110001110110001011110111000;
   assign mem[4605] = 32'b11111110111110001011010101000000;
   assign mem[4606] = 32'b00001001111101000011011000010000;
   assign mem[4607] = 32'b00000110101001011111100011011000;
   assign mem[4608] = 32'b00000100101000011000011101001000;
   assign mem[4609] = 32'b11111010001110010110000111001000;
   assign mem[4610] = 32'b00000111001010111010111001001000;
   assign mem[4611] = 32'b00000101000100111100111110010000;
   assign mem[4612] = 32'b00001000111001010100101010110000;
   assign mem[4613] = 32'b11111011010011011001001010001000;
   assign mem[4614] = 32'b11111100000100111001001111110000;
   assign mem[4615] = 32'b11111111111100000111111010110011;
   assign mem[4616] = 32'b00000000111101110001010000111000;
   assign mem[4617] = 32'b00000011110111111000111111000100;
   assign mem[4618] = 32'b00000001111000110110100000110010;
   assign mem[4619] = 32'b11110110011100111011111011110000;
   assign mem[4620] = 32'b11111011101101010110111100110000;
   assign mem[4621] = 32'b11111010011010100110011100001000;
   assign mem[4622] = 32'b11111011111011111111111010000000;
   assign mem[4623] = 32'b11111010001000010110100100110000;
   assign mem[4624] = 32'b11111110100010010100011111101100;
   assign mem[4625] = 32'b11111111100011001011110111010010;
   assign mem[4626] = 32'b11111110010101000101100010100000;
   assign mem[4627] = 32'b11110110111010111110111110000000;
   assign mem[4628] = 32'b00000100011110100110100110111000;
   assign mem[4629] = 32'b00000111111111001001110101000000;
   assign mem[4630] = 32'b11111101100101110111011001111100;
   assign mem[4631] = 32'b00000011001010101010010110100000;
   assign mem[4632] = 32'b11111111001011000011101111111011;
   assign mem[4633] = 32'b00000000001101111100110110111100;
   assign mem[4634] = 32'b11111110111000011001110101010100;
   assign mem[4635] = 32'b11111101000110011110101100110000;
   assign mem[4636] = 32'b00001000100111011001110011010000;
   assign mem[4637] = 32'b11111110001011100011101001001010;
   assign mem[4638] = 32'b11111100011010010100011000001100;
   assign mem[4639] = 32'b11111111111000110000100010110110;
   assign mem[4640] = 32'b11111110111000111001111100011110;
   assign mem[4641] = 32'b11111100111100011101001000110100;
   assign mem[4642] = 32'b00001000010011111011101001010000;
   assign mem[4643] = 32'b11111111100111110101011011000010;
   assign mem[4644] = 32'b11111010100001001111110111011000;
   assign mem[4645] = 32'b00000100011000000000100110101000;
   assign mem[4646] = 32'b11111001110010101010011101110000;
   assign mem[4647] = 32'b00000100110100110001011100001000;
   assign mem[4648] = 32'b11111101100110001110011101100100;
   assign mem[4649] = 32'b11111100100111101101111100000000;
   assign mem[4650] = 32'b00000001010011000110100001010100;
   assign mem[4651] = 32'b00000010010010100101001111010000;
   assign mem[4652] = 32'b11111101101101100010011011010000;
   assign mem[4653] = 32'b00000010111000011110111101111100;
   assign mem[4654] = 32'b11110100000111001000000010010000;
   assign mem[4655] = 32'b11111110100001001111110110010110;
   assign mem[4656] = 32'b11101100010100101110100010100000;
   assign mem[4657] = 32'b00000011110011101100001100000000;
   assign mem[4658] = 32'b00000101010111011100000110110000;
   assign mem[4659] = 32'b00000010101010101101100010101000;
   assign mem[4660] = 32'b11111110100110111111011101001000;
   assign mem[4661] = 32'b00010111010011000101000000100000;
   assign mem[4662] = 32'b00000100000100011001100001000000;
   assign mem[4663] = 32'b11110001000000101000011001110000;
   assign mem[4664] = 32'b11110000000000011001010001000000;
   assign mem[4665] = 32'b00001101000110010010001111000000;
   assign mem[4666] = 32'b11111100110111101100001010101000;
   assign mem[4667] = 32'b00000101100010000011101110011000;
   assign mem[4668] = 32'b00000010011001101010110111010100;
   assign mem[4669] = 32'b00000001000111100011001011000010;
   assign mem[4670] = 32'b11111110010001000010011001011010;
   assign mem[4671] = 32'b00000011000000011101101101010100;
   assign mem[4672] = 32'b11111011100101110000100110100000;
   assign mem[4673] = 32'b00000101101101011111011001101000;
   assign mem[4674] = 32'b11111111100010010110001010101011;
   assign mem[4675] = 32'b11111110101010000001101011111000;
   assign mem[4676] = 32'b11111100011011000011010011111100;
   assign mem[4677] = 32'b11110110100010110000111000100000;
   assign mem[4678] = 32'b00000010001111000010111010011000;
   assign mem[4679] = 32'b00000011010011000001000111100000;
   assign mem[4680] = 32'b11111010110001100110110010110000;
   assign mem[4681] = 32'b00000000100000011110111010010100;
   assign mem[4682] = 32'b11111100101101010111010100010100;
   assign mem[4683] = 32'b11110111101001100000100111000000;
   assign mem[4684] = 32'b00000001101100000010010000111110;
   assign mem[4685] = 32'b00000101111101101010010010000000;
   assign mem[4686] = 32'b11111101010110010010010011011000;
   assign mem[4687] = 32'b00000101010011000101100100110000;
   assign mem[4688] = 32'b00000000001000011100010010110101;
   assign mem[4689] = 32'b11111110011111001001010110110110;
   assign mem[4690] = 32'b11111001010000000001000101011000;
   assign mem[4691] = 32'b00000100100111000100001001100000;
   assign mem[4692] = 32'b11111010011101101010110011101000;
   assign mem[4693] = 32'b00000000111000011101000011111110;
   assign mem[4694] = 32'b00000000010100101001100111110100;
   assign mem[4695] = 32'b00000001110111110110101100011100;
   assign mem[4696] = 32'b00000001001110000001110111001110;
   assign mem[4697] = 32'b00000000001110011000111110011101;
   assign mem[4698] = 32'b11111101101000010111001110111000;
   assign mem[4699] = 32'b11111111101111110010000110000010;
   assign mem[4700] = 32'b00000001011011111110101011001010;
   assign mem[4701] = 32'b11111111011101010011011001011010;
   assign mem[4702] = 32'b11111110011010101111010010001100;
   assign mem[4703] = 32'b00000010101101110010000011101100;
   assign mem[4704] = 32'b00000010100001000011111001110000;
   assign mem[4705] = 32'b11111011101101011000000110111000;
   assign mem[4706] = 32'b00000000000110010011100110001000;
   assign mem[4707] = 32'b11111000110000011111011001010000;
   assign mem[4708] = 32'b11111111100111001001101110111011;
   assign mem[4709] = 32'b00000011000001001001011000000100;
   assign mem[4710] = 32'b11111110000000010100000110111010;
   assign mem[4711] = 32'b00000010100111011101010011000100;
   assign mem[4712] = 32'b00000001111100000010000100110110;
   assign mem[4713] = 32'b11111001100101111110011001100000;
   assign mem[4714] = 32'b11111110001111001010010010110100;
   assign mem[4715] = 32'b00000000111101101000001011111011;
   assign mem[4716] = 32'b11101011110011001101100110000000;
   assign mem[4717] = 32'b11111011100011011000100100110000;
   assign mem[4718] = 32'b00001100101100100101010110100000;
   assign mem[4719] = 32'b00000101100010100000000010011000;
   assign mem[4720] = 32'b11111011100111000011101000100000;
   assign mem[4721] = 32'b11111110110010101011101011110110;
   assign mem[4722] = 32'b11111101010010010111100110110100;
   assign mem[4723] = 32'b11110110100010001111110000100000;
   assign mem[4724] = 32'b00000011100000111101111110110000;
   assign mem[4725] = 32'b11111111110011000111001011101101;
   assign mem[4726] = 32'b11101101001101001111100100000000;
   assign mem[4727] = 32'b11111001101011000001010111110000;
   assign mem[4728] = 32'b00001001111011011010111010010000;
   assign mem[4729] = 32'b00000101010010001100110100101000;
   assign mem[4730] = 32'b11111111110110000010010010001000;
   assign mem[4731] = 32'b00001011111101011011100110010000;
   assign mem[4732] = 32'b00000000111111110100010011000100;
   assign mem[4733] = 32'b11111101011000001000101101010000;
   assign mem[4734] = 32'b00000110100101111010011010010000;
   assign mem[4735] = 32'b00000001010110110001101100001100;
   assign mem[4736] = 32'b00000101110111001011111000010000;
   assign mem[4737] = 32'b11111111010111110101010110111101;
   assign mem[4738] = 32'b11110111001010100000101010000000;
   assign mem[4739] = 32'b11111011011001000110001011100000;
   assign mem[4740] = 32'b00000000001011101001111101101000;
   assign mem[4741] = 32'b11110110111000101011001000100000;
   assign mem[4742] = 32'b00000101000100101110010100001000;
   assign mem[4743] = 32'b11101101110100101000011011100000;
   assign mem[4744] = 32'b00000110110001010111110011101000;
   assign mem[4745] = 32'b00000000000001111000110011001110;
   assign mem[4746] = 32'b00000010101000010001000111110100;
   assign mem[4747] = 32'b11111111001110111011110000101010;
   assign mem[4748] = 32'b11111110001110111001100110010000;
   assign mem[4749] = 32'b11111110000010111100010101100110;
   assign mem[4750] = 32'b00000110100001010001101101010000;
   assign mem[4751] = 32'b00000011101100011011110011011100;
   assign mem[4752] = 32'b11111101101010100011111111100000;
   assign mem[4753] = 32'b11101111100011110110001110100000;
   assign mem[4754] = 32'b11111101110000010010010101010000;
   assign mem[4755] = 32'b00001000010000111001000010010000;
   assign mem[4756] = 32'b00001001010001010101000110100000;
   assign mem[4757] = 32'b11111100010001010101011001011000;
   assign mem[4758] = 32'b11110111001110001100100000100000;
   assign mem[4759] = 32'b11111111101001001101000001010100;
   assign mem[4760] = 32'b11111110001100101011110111101000;
   assign mem[4761] = 32'b11111100111101100011101001111000;
   assign mem[4762] = 32'b11111100110111111011100010001000;
   assign mem[4763] = 32'b00000101101011010001011010011000;
   assign mem[4764] = 32'b00000001101010010000011010101110;
   assign mem[4765] = 32'b11111110010000011000001010011110;
   assign mem[4766] = 32'b11111101110101100110110010110100;
   assign mem[4767] = 32'b11111110000110001001111100011010;
   assign mem[4768] = 32'b00000000100101101111100011000110;
   assign mem[4769] = 32'b00001010000000111110011010100000;
   assign mem[4770] = 32'b00000110110100110011011110100000;
   assign mem[4771] = 32'b11111000000000110100110100101000;
   assign mem[4772] = 32'b00000011001101100001100000110100;
   assign mem[4773] = 32'b00000000010100110000100111001001;
   assign mem[4774] = 32'b11110101001001101001000100000000;
   assign mem[4775] = 32'b11111110000000000011110011001000;
   assign mem[4776] = 32'b11101110010011001011011000100000;
   assign mem[4777] = 32'b00001010001100100100000010110000;
   assign mem[4778] = 32'b00000010001100111110011001110100;
   assign mem[4779] = 32'b00000110000101000101000010001000;
   assign mem[4780] = 32'b11111011010001010001000100010000;
   assign mem[4781] = 32'b00000011010101010001101011000000;
   assign mem[4782] = 32'b11111111100011111001001001011100;
   assign mem[4783] = 32'b11110110111000001010110000100000;
   assign mem[4784] = 32'b00000010111100010100110101111100;
   assign mem[4785] = 32'b00000011011111010001110110011100;
   assign mem[4786] = 32'b00000100010111011101100010111000;
   assign mem[4787] = 32'b00000010001010111101000100101100;
   assign mem[4788] = 32'b11110111011101001001110110010000;
   assign mem[4789] = 32'b11111000110010000100000010111000;
   assign mem[4790] = 32'b11111100011011111011001000111100;
   assign mem[4791] = 32'b00000011011001000000000110100100;
   assign mem[4792] = 32'b00000100011111100010010010111000;
   assign mem[4793] = 32'b11111111011100001110000011000011;
   assign mem[4794] = 32'b11111001001000010010010110100000;
   assign mem[4795] = 32'b00000100011011011010110111111000;
   assign mem[4796] = 32'b11110111001011011100000101010000;
   assign mem[4797] = 32'b00000011100100010101101010011000;
   assign mem[4798] = 32'b11111101010010000000111011010000;
   assign mem[4799] = 32'b11111011101011111110010110010000;
   assign mem[4800] = 32'b00000000110011001101000101101010;
   assign mem[4801] = 32'b00000000011001001011000101101100;
   assign mem[4802] = 32'b11111111001111011101110100001100;
   assign mem[4803] = 32'b11111011100110001110010011101000;
   assign mem[4804] = 32'b00000010011001110010011111101000;
   assign mem[4805] = 32'b11111111010010001111000101110010;
   assign mem[4806] = 32'b11111111011110101111100111011110;
   assign mem[4807] = 32'b11111110001110111000111001001010;
   assign mem[4808] = 32'b11111101111111011111010101111000;
   assign mem[4809] = 32'b00000000111010110100101011111100;
   assign mem[4810] = 32'b00000001001010010010001010111110;
   assign mem[4811] = 32'b11111101010111110011111000011100;
   assign mem[4812] = 32'b11111101000000011100110111101000;
   assign mem[4813] = 32'b11110001011010010010101100000000;
   assign mem[4814] = 32'b00000000001110111010011010100110;
   assign mem[4815] = 32'b00000101001101101001110101010000;
   assign mem[4816] = 32'b00000011110101000001000010100100;
   assign mem[4817] = 32'b11111101011100010001010011000000;
   assign mem[4818] = 32'b11111011011101011010100110001000;
   assign mem[4819] = 32'b00000000011100000101000110001010;
   assign mem[4820] = 32'b00000011000000110011100101111000;
   assign mem[4821] = 32'b11110110010100111111011111010000;
   assign mem[4822] = 32'b00000010010010101111100101011000;
   assign mem[4823] = 32'b11111100111101011001011010110000;
   assign mem[4824] = 32'b11110100001101011110100011000000;
   assign mem[4825] = 32'b00000010110001101011111010001000;
   assign mem[4826] = 32'b11111100000100101101011100111000;
   assign mem[4827] = 32'b00000110101100111101010100000000;
   assign mem[4828] = 32'b00000000010100111000111110010001;
   assign mem[4829] = 32'b00000000010011101110101000001010;
   assign mem[4830] = 32'b00000010011100011101101101101000;
   assign mem[4831] = 32'b00001100101110011111111010100000;
   assign mem[4832] = 32'b00001001000001010001110010000000;
   assign mem[4833] = 32'b11111101000010001011000110011000;
   assign mem[4834] = 32'b00000101001101010001011010101000;
   assign mem[4835] = 32'b00000000010011110001000101110011;
   assign mem[4836] = 32'b00001000010010100101011000100000;
   assign mem[4837] = 32'b11101000100000011000010100000000;
   assign mem[4838] = 32'b11110111110100100111110111010000;
   assign mem[4839] = 32'b11111010010110010100000100010000;
   assign mem[4840] = 32'b11111110110001010100001010110110;
   assign mem[4841] = 32'b11111011000111010110000101110000;
   assign mem[4842] = 32'b00000010110111010110110100111000;
   assign mem[4843] = 32'b11111001101000011100101100011000;
   assign mem[4844] = 32'b11111001101101001111001000101000;
   assign mem[4845] = 32'b00000101100000110011111100000000;
   assign mem[4846] = 32'b00000010010010011000111111101000;
   assign mem[4847] = 32'b00000011101001101000001100110000;
   assign mem[4848] = 32'b00000010110011101110100011001000;
   assign mem[4849] = 32'b11110100001110100001111000100000;
   assign mem[4850] = 32'b00000010010110111110110110011000;
   assign mem[4851] = 32'b11111000111000011011000011101000;
   assign mem[4852] = 32'b11111111000000111110000011101111;
   assign mem[4853] = 32'b11111110000000111110100110100100;
   assign mem[4854] = 32'b11110110100010101011101010100000;
   assign mem[4855] = 32'b11111110000010010101110100010100;
   assign mem[4856] = 32'b11110110100010011111110100000000;
   assign mem[4857] = 32'b00000011010001111001111111011100;
   assign mem[4858] = 32'b00000101111000110111111111111000;
   assign mem[4859] = 32'b00001001011100000111101011000000;
   assign mem[4860] = 32'b11111110011111110101111101101110;
   assign mem[4861] = 32'b00000100000000000001110110011000;
   assign mem[4862] = 32'b11111111000101011111111111001000;
   assign mem[4863] = 32'b11111001001100111001111110100000;
   assign mem[4864] = 32'b00000011011000101001010100110100;
   assign mem[4865] = 32'b00000111000000101100111110100000;
   assign mem[4866] = 32'b11111101111111000110010101111100;
   assign mem[4867] = 32'b00000100010111110001000001001000;
   assign mem[4868] = 32'b11111100101110100100000011000100;
   assign mem[4869] = 32'b00000101010001010011010001011000;
   assign mem[4870] = 32'b11111011100001001110100100111000;
   assign mem[4871] = 32'b00000101101000010000101011100000;
   assign mem[4872] = 32'b00000000110010111100110111110000;
   assign mem[4873] = 32'b00001001000111110110000001010000;
   assign mem[4874] = 32'b11110101010110011010001000100000;
   assign mem[4875] = 32'b11111000011111001001000110001000;
   assign mem[4876] = 32'b11111010001011000101111011010000;
   assign mem[4877] = 32'b00001000111010010011101110000000;
   assign mem[4878] = 32'b11101110011100111000001000000000;
   assign mem[4879] = 32'b11110101001110100111000010100000;
   assign mem[4880] = 32'b00000110001100111101110000100000;
   assign mem[4881] = 32'b11111100011101110100111101100000;
   assign mem[4882] = 32'b00000101110010001101100110001000;
   assign mem[4883] = 32'b11111000011111110001110100110000;
   assign mem[4884] = 32'b11110000011110011101001111000000;
   assign mem[4885] = 32'b00000001100100000000011000101010;
   assign mem[4886] = 32'b11111001010111111100011101011000;
   assign mem[4887] = 32'b00000100011110010111110110010000;
   assign mem[4888] = 32'b00001000110100001011001100000000;
   assign mem[4889] = 32'b00000001011111011111111000000000;
   assign mem[4890] = 32'b11110110001111001110111000110000;
   assign mem[4891] = 32'b11111110011101110000010110000100;
   assign mem[4892] = 32'b00000010111010111101110101011100;
   assign mem[4893] = 32'b00000000001011101101101001101100;
   assign mem[4894] = 32'b11111110111011000011010101001000;
   assign mem[4895] = 32'b00000011000010010111101100001100;
   assign mem[4896] = 32'b00000011100111000010101010001100;
   assign mem[4897] = 32'b00000110110010111001100100100000;
   assign mem[4898] = 32'b11111100101011100010010100110000;
   assign mem[4899] = 32'b11111100010010110110100011001000;
   assign mem[4900] = 32'b11111111100010100110010110000101;
   assign mem[4901] = 32'b00000100000100000100101001110000;
   assign mem[4902] = 32'b00000100100000000101010111110000;
   assign mem[4903] = 32'b00000011111110111011110111010000;
   assign mem[4904] = 32'b11110000011111111101001000000000;
   assign mem[4905] = 32'b11110111010100001000000011110000;
   assign mem[4906] = 32'b11111101111010101101110101110000;
   assign mem[4907] = 32'b00000110100001010100111001110000;
   assign mem[4908] = 32'b11110011101000001010111101010000;
   assign mem[4909] = 32'b11111001101100110000111111001000;
   assign mem[4910] = 32'b11110110110100100011110100110000;
   assign mem[4911] = 32'b00000001110000100111011010011010;
   assign mem[4912] = 32'b00000110100000101000111000001000;
   assign mem[4913] = 32'b00000010110010110101010100000000;
   assign mem[4914] = 32'b00001011100101101100011010000000;
   assign mem[4915] = 32'b11111011001001001000101111011000;
   assign mem[4916] = 32'b11111100000110001011010110001100;
   assign mem[4917] = 32'b00000101100000100010101111010000;
   assign mem[4918] = 32'b11110101000010111110111011100000;
   assign mem[4919] = 32'b11110001111010011000000110000000;
   assign mem[4920] = 32'b11111100010001010001000000010100;
   assign mem[4921] = 32'b00000010000000011011111010010100;
   assign mem[4922] = 32'b11111100101110100100111101110100;
   assign mem[4923] = 32'b11111011000100100010100101000000;
   assign mem[4924] = 32'b11111110000111101100110010010110;
   assign mem[4925] = 32'b00001000001000111100111010010000;
   assign mem[4926] = 32'b00000011001110001111101100001100;
   assign mem[4927] = 32'b11110101100110011000011111110000;
   assign mem[4928] = 32'b11111110010101110000110001111110;
   assign mem[4929] = 32'b00000101010100001011101101000000;
   assign mem[4930] = 32'b00000010011001111110110000111000;
   assign mem[4931] = 32'b00000000010101101100010110101000;
   assign mem[4932] = 32'b00000111000010000001011100001000;
   assign mem[4933] = 32'b11111111000111010000110010111010;
   assign mem[4934] = 32'b11110110110000001100011000010000;
   assign mem[4935] = 32'b11111001110011010001011001101000;
   assign mem[4936] = 32'b11111000100111101110011100110000;
   assign mem[4937] = 32'b00000101100110100011010101100000;
   assign mem[4938] = 32'b11111101010100000101001000110100;
   assign mem[4939] = 32'b00000110001010111100100100010000;
   assign mem[4940] = 32'b11110001110110011010001010010000;
   assign mem[4941] = 32'b00000010110110010111100110010100;
   assign mem[4942] = 32'b00000100000110111100001101011000;
   assign mem[4943] = 32'b00000001011001011110001000001100;
   assign mem[4944] = 32'b11111100001111100101100111001000;
   assign mem[4945] = 32'b11110111011001011000111110110000;
   assign mem[4946] = 32'b11111000001101010011100101110000;
   assign mem[4947] = 32'b00000111101011010001010001011000;
   assign mem[4948] = 32'b00000010111000101100001101110000;
   assign mem[4949] = 32'b11111100011111111000010111010100;
   assign mem[4950] = 32'b11111011101101000100110100001000;
   assign mem[4951] = 32'b11111111000011111000000000111000;
   assign mem[4952] = 32'b11111110111000000100011111101000;
   assign mem[4953] = 32'b11111101101100111101110111111000;
   assign mem[4954] = 32'b11111101011110101010101100100100;
   assign mem[4955] = 32'b00000010001001001110111100111100;
   assign mem[4956] = 32'b00000001010010111011010100101010;
   assign mem[4957] = 32'b00000001100000100101001110010100;
   assign mem[4958] = 32'b00000000100011000000101111110000;
   assign mem[4959] = 32'b00000000010000100111101010110001;
   assign mem[4960] = 32'b00000111000101111011100000101000;
   assign mem[4961] = 32'b11111010010011101010011000101000;
   assign mem[4962] = 32'b00000010111001010101000111100000;
   assign mem[4963] = 32'b00000010001110101001001000001000;
   assign mem[4964] = 32'b11110010110101100100001001100000;
   assign mem[4965] = 32'b00000001110010110001110100001110;
   assign mem[4966] = 32'b11111100111011001011111110101000;
   assign mem[4967] = 32'b00000100000111001001000111100000;
   assign mem[4968] = 32'b00000000010101111010000000100111;
   assign mem[4969] = 32'b11111110000101101001011111010100;
   assign mem[4970] = 32'b00000010100101001111001001111100;
   assign mem[4971] = 32'b00000011001110001111010010000100;
   assign mem[4972] = 32'b11111111110000111100010101010111;
   assign mem[4973] = 32'b11110001011110111101011111100000;
   assign mem[4974] = 32'b11111101101111101000010101100000;
   assign mem[4975] = 32'b00000000101010000001111001100100;
   assign mem[4976] = 32'b00000011110011010010110010110000;
   assign mem[4977] = 32'b11111110010101101111110001010000;
   assign mem[4978] = 32'b11111001010110000011010101000000;
   assign mem[4979] = 32'b00000010010011110011011001111100;
   assign mem[4980] = 32'b00000001001011000000101000011010;
   assign mem[4981] = 32'b11111111000001100111100100111110;
   assign mem[4982] = 32'b11111000011000001011101100111000;
   assign mem[4983] = 32'b00000010001000011000011100101100;
   assign mem[4984] = 32'b00000010000100000100111111010000;
   assign mem[4985] = 32'b11111100000111111110011101111000;
   assign mem[4986] = 32'b00001001001100111000010111100000;
   assign mem[4987] = 32'b11111010001010101111011010000000;
   assign mem[4988] = 32'b11111101000010011000010101101100;
   assign mem[4989] = 32'b00000100010011101011111110011000;
   assign mem[4990] = 32'b11110011111001110001110001100000;
   assign mem[4991] = 32'b00000111101110001010111000101000;
   assign mem[4992] = 32'b00000110011000011111111101100000;
   assign mem[4993] = 32'b11111101111001011111011101010100;
   assign mem[4994] = 32'b11111101111100001011011111110100;
   assign mem[4995] = 32'b11111001011000110001111000101000;
   assign mem[4996] = 32'b11111101010000011101001001111000;
   assign mem[4997] = 32'b11111110101100100111110000100000;
   assign mem[4998] = 32'b11111111011010110101010111001110;
   assign mem[4999] = 32'b11110011001001100100110011100000;
   assign mem[5000] = 32'b11111101000011100011101101110000;
   assign mem[5001] = 32'b11111010011101000101100110110000;
   assign mem[5002] = 32'b00000000111111000011100100001110;
   assign mem[5003] = 32'b00000001101000110010110101001110;
   assign mem[5004] = 32'b11110100101011000011100001110000;
   assign mem[5005] = 32'b11111110010010010111101111001110;
   assign mem[5006] = 32'b11111010101100100011001001010000;
   assign mem[5007] = 32'b00000001101011111011110110111100;
   assign mem[5008] = 32'b11111111000001001011010000110110;
   assign mem[5009] = 32'b00000011011010011000111011111000;
   assign mem[5010] = 32'b11111000001000010111111001101000;
   assign mem[5011] = 32'b11110100000011101110110000100000;
   assign mem[5012] = 32'b00000000110011000011000010101100;
   assign mem[5013] = 32'b00000000100101001011011110011100;
   assign mem[5014] = 32'b11110100101101110101010011010000;
   assign mem[5015] = 32'b00000010101000101100010100111100;
   assign mem[5016] = 32'b11111101111100000010010010011100;
   assign mem[5017] = 32'b00000011001111010011111100110100;
   assign mem[5018] = 32'b00000000001000100000101110011110;
   assign mem[5019] = 32'b00000110110011111100011110001000;
   assign mem[5020] = 32'b11111111000000110010000111001101;
   assign mem[5021] = 32'b11111110110001001010111110100000;
   assign mem[5022] = 32'b00000111000111011100110011110000;
   assign mem[5023] = 32'b00000000011001000100100101110011;
   assign mem[5024] = 32'b11111001011000000110101001000000;
   assign mem[5025] = 32'b11111111101010001000110010011111;
   assign mem[5026] = 32'b11111110001100011100101010010100;
   assign mem[5027] = 32'b00000010011001000101010000000100;
   assign mem[5028] = 32'b11111100011100111101111000000000;
   assign mem[5029] = 32'b11111011111000011111100111100000;
   assign mem[5030] = 32'b11111101110101010101001000011000;
   assign mem[5031] = 32'b00000001010110110110011110101110;
   assign mem[5032] = 32'b00000010110101100000100010001000;
   assign mem[5033] = 32'b11111100011111011111010000001000;
   assign mem[5034] = 32'b00000111111010100010101111010000;
   assign mem[5035] = 32'b11111101001001000110111011100000;
   assign mem[5036] = 32'b00000010100111010000010100011100;
   assign mem[5037] = 32'b11111010010011110101101110111000;
   assign mem[5038] = 32'b00000001110100011111011111101110;
   assign mem[5039] = 32'b00000010101010000100110001010100;
   assign mem[5040] = 32'b00000100011101101000011110110000;
   assign mem[5041] = 32'b00000111011010111000100100001000;
   assign mem[5042] = 32'b00000010100000000000010000110000;
   assign mem[5043] = 32'b00000011000000110111001110111100;
   assign mem[5044] = 32'b00001000101100001000000111000000;
   assign mem[5045] = 32'b11111110001001100101010111011000;
   assign mem[5046] = 32'b11111101101100000011000100110000;
   assign mem[5047] = 32'b00000000100100100010101001001010;
   assign mem[5048] = 32'b00000000000110100101110100111001;
   assign mem[5049] = 32'b11110000111010111000001001100000;
   assign mem[5050] = 32'b11111101100010011100000101010000;
   assign mem[5051] = 32'b11111111101101111001101010110100;
   assign mem[5052] = 32'b00000101111011101100011001010000;
   assign mem[5053] = 32'b00000101011010010010111010110000;
   assign mem[5054] = 32'b11110010111011001001101011000000;
   assign mem[5055] = 32'b11111100111011001100100011010100;
   assign mem[5056] = 32'b11110111010011001000111100000000;
   assign mem[5057] = 32'b00000011100110100011101011111000;
   assign mem[5058] = 32'b00000011100010001101100100110100;
   assign mem[5059] = 32'b11111111011101011010111101010000;
   assign mem[5060] = 32'b00000101100110110110100111110000;
   assign mem[5061] = 32'b11111101001100111111111001101100;
   assign mem[5062] = 32'b00000011100101100011010100011100;
   assign mem[5063] = 32'b11111101000010111011000110010000;
   assign mem[5064] = 32'b00000011000110011001111100101100;
   assign mem[5065] = 32'b11111110100000001011111000001010;
   assign mem[5066] = 32'b11111110101111100000011101110010;
   assign mem[5067] = 32'b00000110001100100001111100010000;
   assign mem[5068] = 32'b11110110000011101000011101110000;
   assign mem[5069] = 32'b11110101000000101011101101010000;
   assign mem[5070] = 32'b00000000000100100101001101010110;
   assign mem[5071] = 32'b11111111101111100010100010011001;
   assign mem[5072] = 32'b00000000010100000110111101011100;
   assign mem[5073] = 32'b11111100011010001001111001001100;
   assign mem[5074] = 32'b00000010010111101001001000001100;
   assign mem[5075] = 32'b11111101001110010000001000010000;
   assign mem[5076] = 32'b11111000000100010111011001011000;
   assign mem[5077] = 32'b00000110011100110000101110111000;
   assign mem[5078] = 32'b11111111100100100001100000111110;
   assign mem[5079] = 32'b00000000000110010001111011010001;
   assign mem[5080] = 32'b00000010101100011010101110100100;
   assign mem[5081] = 32'b00000011000010100101110111011000;
   assign mem[5082] = 32'b11111101010000010010110100111000;
   assign mem[5083] = 32'b00000100011111011111100001001000;
   assign mem[5084] = 32'b11111110010110010001000111111100;
   assign mem[5085] = 32'b11111110000000111111010110101000;
   assign mem[5086] = 32'b00000100001101011100010100110000;
   assign mem[5087] = 32'b00000000111011000111000000101110;
   assign mem[5088] = 32'b11111000111000001001001110100000;
   assign mem[5089] = 32'b00000010000101101000101100110000;
   assign mem[5090] = 32'b00000110111111101100011010010000;
   assign mem[5091] = 32'b00000001100100000000110101010000;
   assign mem[5092] = 32'b00000000001000101001100000001100;
   assign mem[5093] = 32'b11101011010101001010010011000000;
   assign mem[5094] = 32'b11111110110001001010000100010000;
   assign mem[5095] = 32'b00000010100001100110011100011100;
   assign mem[5096] = 32'b00000100111110111010001101110000;
   assign mem[5097] = 32'b11111010100111010011010101100000;
   assign mem[5098] = 32'b11111101011100001000100000110000;
   assign mem[5099] = 32'b11111101010110100011111110011000;
   assign mem[5100] = 32'b11111011011101001100000111110000;
   assign mem[5101] = 32'b00000100101000001001100100101000;
   assign mem[5102] = 32'b00000010100101010111101111010100;
   assign mem[5103] = 32'b11110110011000100000010000010000;
   assign mem[5104] = 32'b00000100000101110111011011000000;
   assign mem[5105] = 32'b00001010101011110000011010010000;
   assign mem[5106] = 32'b00000001000010001011011111110010;
   assign mem[5107] = 32'b11110100110001000110110101100000;
   assign mem[5108] = 32'b00000000110111001000110001001011;
   assign mem[5109] = 32'b11110101010010000110000010110000;
   assign mem[5110] = 32'b11110101000011100001101010110000;
   assign mem[5111] = 32'b00000010110100000100111001010000;
   assign mem[5112] = 32'b00000001010001111000110011111110;
   assign mem[5113] = 32'b11110110100001011100001100000000;
   assign mem[5114] = 32'b00000001000011110000100111111100;
   assign mem[5115] = 32'b00000101111110000100000100110000;
   assign mem[5116] = 32'b00000001000110110001011011100010;
   assign mem[5117] = 32'b11111110000011010100010100110100;
   assign mem[5118] = 32'b11111100001100011100000100011100;
   assign mem[5119] = 32'b11111011111000100101011101101000;
   assign mem[5120] = 32'b11111011111001101100010010010000;
   assign mem[5121] = 32'b11110011010100011010001111100000;
   assign mem[5122] = 32'b11111011110110001100010011110000;
   assign mem[5123] = 32'b00000101111011010111000001100000;
   assign mem[5124] = 32'b11110100000111111111110111010000;
   assign mem[5125] = 32'b00000000011010010000000011110010;
   assign mem[5126] = 32'b00000011101000110100111111110100;
   assign mem[5127] = 32'b11110101011101011111111011100000;
   assign mem[5128] = 32'b00000111000110110010010010100000;
   assign mem[5129] = 32'b00000101001000100111001111000000;
   assign mem[5130] = 32'b00000111011100101001001001011000;
   assign mem[5131] = 32'b00000001111100011010110001100110;
   assign mem[5132] = 32'b00000100010100000101010100110000;
   assign mem[5133] = 32'b00000101100000010010010010011000;
   assign mem[5134] = 32'b11111011111000100010111000000000;
   assign mem[5135] = 32'b11101101010100001100001001000000;
   assign mem[5136] = 32'b11110101101111101111111001110000;
   assign mem[5137] = 32'b11111110101000010011110001111010;
   assign mem[5138] = 32'b11111001111010111011001100001000;
   assign mem[5139] = 32'b00000011000100101100001100111100;
   assign mem[5140] = 32'b00000100001010101101010101000000;
   assign mem[5141] = 32'b11111101011100101010001001101000;
   assign mem[5142] = 32'b00000001011100110110101001010100;
   assign mem[5143] = 32'b11111101110100111110110010101100;
   assign mem[5144] = 32'b11110110000000100101111010010000;
   assign mem[5145] = 32'b00000000110001000010001010010010;
   assign mem[5146] = 32'b11111010101111001110010100010000;
   assign mem[5147] = 32'b11111111110111010011111001010010;
   assign mem[5148] = 32'b11111110111011011001101010101000;
   assign mem[5149] = 32'b11111110010110000011001111101100;
   assign mem[5150] = 32'b11111011010011111000000011001000;
   assign mem[5151] = 32'b11110000101110000101110110110000;
   assign mem[5152] = 32'b11111011111110000101000011100000;
   assign mem[5153] = 32'b00000010011000010000010000110100;
   assign mem[5154] = 32'b11110101001011000111100111100000;
   assign mem[5155] = 32'b00000110101011011111000010000000;
   assign mem[5156] = 32'b11111100010001011111010000110100;
   assign mem[5157] = 32'b00000111000000000000010111001000;
   assign mem[5158] = 32'b11111110101111010101001011010000;
   assign mem[5159] = 32'b00000100000000010111010010100000;
   assign mem[5160] = 32'b11111101110111011101001000110100;
   assign mem[5161] = 32'b11111110010100001001011000001100;
   assign mem[5162] = 32'b11111111001001111100100100101001;
   assign mem[5163] = 32'b11110011010001110111100100000000;
   assign mem[5164] = 32'b11111011101011111110010011111000;
   assign mem[5165] = 32'b00001100110100011101100100010000;
   assign mem[5166] = 32'b00000110110100100000010100110000;
   assign mem[5167] = 32'b11111010010001111011010101010000;
   assign mem[5168] = 32'b11111001110011101100111010100000;
   assign mem[5169] = 32'b00000010110110011011110110110000;
   assign mem[5170] = 32'b11111100010101110001010000110000;
   assign mem[5171] = 32'b00000010000110011111001001011000;
   assign mem[5172] = 32'b00000001100110001110111101000100;
   assign mem[5173] = 32'b11111111100100010100011100010101;
   assign mem[5174] = 32'b00000101000000111000010111100000;
   assign mem[5175] = 32'b11111001110111101001111000111000;
   assign mem[5176] = 32'b00000101000000010001110001010000;
   assign mem[5177] = 32'b11111010000110011001011111010000;
   assign mem[5178] = 32'b11111101101110011111111001111000;
   assign mem[5179] = 32'b00000001011000001010100100001000;
   assign mem[5180] = 32'b11110101101101011111110101000000;
   assign mem[5181] = 32'b00000101011011010010101111011000;
   assign mem[5182] = 32'b11111111110100111000011010001000;
   assign mem[5183] = 32'b00000000001010010101001110110010;
   assign mem[5184] = 32'b00000001000111011011101101011110;
   assign mem[5185] = 32'b11111100110101010110101110101000;
   assign mem[5186] = 32'b00000001001100000101100011111100;
   assign mem[5187] = 32'b00000010011101100000010100001100;
   assign mem[5188] = 32'b11111101110010101001110110011100;
   assign mem[5189] = 32'b00000011110101010000000100010000;
   assign mem[5190] = 32'b11111110101001110100000110101000;
   assign mem[5191] = 32'b11111111111011110101110111011000;
   assign mem[5192] = 32'b00000000001000101000001110001101;
   assign mem[5193] = 32'b11111111110101100111100010110110;
   assign mem[5194] = 32'b00000010100110000010110111010100;
   assign mem[5195] = 32'b11111110010111100010100111011110;
   assign mem[5196] = 32'b00000011011110110110010011011000;
   assign mem[5197] = 32'b00000011000011111101001011111100;
   assign mem[5198] = 32'b11111110001001000100011110100100;
   assign mem[5199] = 32'b11111101101110100010011111110000;
   assign mem[5200] = 32'b00000010101110001011111011011100;
   assign mem[5201] = 32'b11111100110101001111011000110100;
   assign mem[5202] = 32'b11111100100111100110100110101000;
   assign mem[5203] = 32'b11111011000110110010110011110000;
   assign mem[5204] = 32'b11110111001010101010001001000000;
   assign mem[5205] = 32'b00000101011100101111001000111000;
   assign mem[5206] = 32'b00000111001000011011110010001000;
   assign mem[5207] = 32'b00000101101110111001011010001000;
   assign mem[5208] = 32'b11110111111001111001100110100000;
   assign mem[5209] = 32'b11111001100101100111010110011000;
   assign mem[5210] = 32'b00000010011110011111001111010000;
   assign mem[5211] = 32'b00000110111101111001111110011000;
   assign mem[5212] = 32'b00001010100001000110001001000000;
   assign mem[5213] = 32'b11110110010111000101011011010000;
   assign mem[5214] = 32'b00000100001100111101001100100000;
   assign mem[5215] = 32'b00000000001001011101010010001111;
   assign mem[5216] = 32'b11111010100101001000000010100000;
   assign mem[5217] = 32'b11110110111101011010101101000000;
   assign mem[5218] = 32'b00000010000111011100001001111000;
   assign mem[5219] = 32'b11111111101011110100110001101100;
   assign mem[5220] = 32'b11111101110011001100100101101000;
   assign mem[5221] = 32'b11111110101100101000111110011110;
   assign mem[5222] = 32'b11111000011110010100110000110000;
   assign mem[5223] = 32'b00000000110001110111100001010001;
   assign mem[5224] = 32'b11110111000110011010001110000000;
   assign mem[5225] = 32'b00000110001100000100000011000000;
   assign mem[5226] = 32'b11111011111011001111111110111000;
   assign mem[5227] = 32'b00000100000110110010101101101000;
   assign mem[5228] = 32'b00000010101111111010111101111100;
   assign mem[5229] = 32'b00000001001111110001010101000100;
   assign mem[5230] = 32'b00000001010100001010011101011000;
   assign mem[5231] = 32'b11111010000001001011100100110000;
   assign mem[5232] = 32'b00000011101110011111001001100100;
   assign mem[5233] = 32'b11111011000010111011110111110000;
   assign mem[5234] = 32'b11111011111011110111110011001000;
   assign mem[5235] = 32'b00000001001100110110111100111010;
   assign mem[5236] = 32'b11111000111010110111111110101000;
   assign mem[5237] = 32'b00000101111000101010000011101000;
   assign mem[5238] = 32'b00000001001111110010100011100100;
   assign mem[5239] = 32'b11111011111010010011010001000000;
   assign mem[5240] = 32'b11111010000111000000111001011000;
   assign mem[5241] = 32'b11110110001110000100111111100000;
   assign mem[5242] = 32'b11110111101100111100001101000000;
   assign mem[5243] = 32'b00001001111110100101111011100000;
   assign mem[5244] = 32'b11111110000001011011001111111100;
   assign mem[5245] = 32'b00000011010100111010101001000000;
   assign mem[5246] = 32'b00000111101101000110111111000000;
   assign mem[5247] = 32'b00000111111001011100100110001000;
   assign mem[5248] = 32'b11111100100111000100110101011000;
   assign mem[5249] = 32'b11101110010100001101110110100000;
   assign mem[5250] = 32'b11111101001100001000111011010100;
   assign mem[5251] = 32'b00000001100011011100100110000110;
   assign mem[5252] = 32'b11111111001001010100000000011111;
   assign mem[5253] = 32'b11111110111110111001110001100100;
   assign mem[5254] = 32'b11111000001101111001110100111000;
   assign mem[5255] = 32'b00000010000000010000010000011000;
   assign mem[5256] = 32'b00000101110000110011001010001000;
   assign mem[5257] = 32'b00000010111010000111100010100000;
   assign mem[5258] = 32'b11111001110011011101001011011000;
   assign mem[5259] = 32'b11111110110101011010000000010010;
   assign mem[5260] = 32'b11111010101001110000100100010000;
   assign mem[5261] = 32'b11111001011111111000101001111000;
   assign mem[5262] = 32'b11110110111101100010101110110000;
   assign mem[5263] = 32'b00001010000011110111001010110000;
   assign mem[5264] = 32'b00000001010000011010001101011010;
   assign mem[5265] = 32'b11111111010110011110110011010110;
   assign mem[5266] = 32'b11111001000111001001111111001000;
   assign mem[5267] = 32'b00000001110001011010000000111010;
   assign mem[5268] = 32'b00000010001111101000110101011000;
   assign mem[5269] = 32'b11111110100101111111100010111000;
   assign mem[5270] = 32'b11111110001110111111101110100000;
   assign mem[5271] = 32'b00000001110101001100000001001000;
   assign mem[5272] = 32'b00000101000110001000001110111000;
   assign mem[5273] = 32'b00000010101110100101100111111000;
   assign mem[5274] = 32'b00000001001110011001010100101100;
   assign mem[5275] = 32'b11101000010100100111101011000000;
   assign mem[5276] = 32'b00000000111000011100011011100101;
   assign mem[5277] = 32'b00000001100000110110100111100100;
   assign mem[5278] = 32'b11111100111001010110011101010000;
   assign mem[5279] = 32'b00000010101100001001001110000100;
   assign mem[5280] = 32'b11111111101001101111111111111001;
   assign mem[5281] = 32'b11111001010101101111100010110000;
   assign mem[5282] = 32'b00000000111010010111111111011001;
   assign mem[5283] = 32'b11111111011010100001000111001001;
   assign mem[5284] = 32'b11111000010111111111111001111000;
   assign mem[5285] = 32'b00001000100100010101100010010000;
   assign mem[5286] = 32'b11111100110101010110111101011100;
   assign mem[5287] = 32'b00000000011001010101010111010011;
   assign mem[5288] = 32'b00000010000100011101001101110000;
   assign mem[5289] = 32'b00000100100101001010101101101000;
   assign mem[5290] = 32'b11111110101111110000100100101100;
   assign mem[5291] = 32'b11111100101111001010000101100100;
   assign mem[5292] = 32'b11111111010001111110111100010000;
   assign mem[5293] = 32'b00000100000111000000010000111000;
   assign mem[5294] = 32'b00000010000010110010001001110000;
   assign mem[5295] = 32'b00000000101000010000110010001101;
   assign mem[5296] = 32'b11110101001100101000110101010000;
   assign mem[5297] = 32'b00001001110000111101111110000000;
   assign mem[5298] = 32'b11111110010100101100000111100000;
   assign mem[5299] = 32'b11111100101100011101001011011000;
   assign mem[5300] = 32'b00000000111111010011100111101101;
   assign mem[5301] = 32'b00000110010111110000111011111000;
   assign mem[5302] = 32'b00000101010111011001010001100000;
   assign mem[5303] = 32'b11111101110011110111010000111000;
   assign mem[5304] = 32'b11110111001111111101101011010000;
   assign mem[5305] = 32'b00001000000011111110001101010000;
   assign mem[5306] = 32'b00001000001110111101101001100000;
   assign mem[5307] = 32'b11111011101000001010110011010000;
   assign mem[5308] = 32'b11110110100011111001011011000000;
   assign mem[5309] = 32'b00000011000111001100000100001100;
   assign mem[5310] = 32'b11101111000001001111101100000000;
   assign mem[5311] = 32'b11101111000110100000100100100000;
   assign mem[5312] = 32'b00000001111111101010101111010000;
   assign mem[5313] = 32'b00000110101111001010111100000000;
   assign mem[5314] = 32'b11110001000011100110111000110000;
   assign mem[5315] = 32'b00000011001011001010101000011000;
   assign mem[5316] = 32'b00000000100111100000000000111100;
   assign mem[5317] = 32'b11111101110001011111000101001100;
   assign mem[5318] = 32'b00001000111100011000110001100000;
   assign mem[5319] = 32'b00000011110010110111011111000000;
   assign mem[5320] = 32'b11111101000111001111110010111000;
   assign mem[5321] = 32'b00001010001000001111011000110000;
   assign mem[5322] = 32'b00000110011010001100100111110000;
   assign mem[5323] = 32'b11111100101110101101110101010100;
   assign mem[5324] = 32'b00000110100011011010100100000000;
   assign mem[5325] = 32'b11110100101110111010000010110000;
   assign mem[5326] = 32'b11110000011000101111000000010000;
   assign mem[5327] = 32'b00000111000010101011100001010000;
   assign mem[5328] = 32'b11111011110011001111100100000000;
   assign mem[5329] = 32'b11111110101001010010100101000010;
   assign mem[5330] = 32'b11111010101100010001110000100000;
   assign mem[5331] = 32'b11111011000111101001101110111000;
   assign mem[5332] = 32'b11111001110011111110100100010000;
   assign mem[5333] = 32'b00000011011010011111000000000100;
   assign mem[5334] = 32'b11110011101001011000100010000000;
   assign mem[5335] = 32'b00000111100000111010010000000000;
   assign mem[5336] = 32'b11111101101010010101101100101100;
   assign mem[5337] = 32'b00000001010011010001100111101010;
   assign mem[5338] = 32'b00000001011110001110111111100010;
   assign mem[5339] = 32'b00000010110011110010010100111100;
   assign mem[5340] = 32'b11111101000110000101100001011000;
   assign mem[5341] = 32'b11111011000010000001011111101000;
   assign mem[5342] = 32'b11111101100101000011010011101100;
   assign mem[5343] = 32'b00001001111000111010111011010000;
   assign mem[5344] = 32'b11111110101000101000111011100010;
   assign mem[5345] = 32'b11111110000111010000000000010110;
   assign mem[5346] = 32'b11111111110111011010010110101011;
   assign mem[5347] = 32'b00000000010000000010110111011011;
   assign mem[5348] = 32'b00000100101100000100010101110000;
   assign mem[5349] = 32'b00000010011011000000110110001000;
   assign mem[5350] = 32'b00001000101011011111000110100000;
   assign mem[5351] = 32'b11111111001010110000101110001010;
   assign mem[5352] = 32'b00000101011111111001110010010000;
   assign mem[5353] = 32'b11111111010001111100110010110011;
   assign mem[5354] = 32'b11111101101101111001100110111000;
   assign mem[5355] = 32'b00000010001101101100001001011100;
   assign mem[5356] = 32'b11101010101001001110001110100000;
   assign mem[5357] = 32'b00000101000101011111001100000000;
   assign mem[5358] = 32'b11111110111010101001111110001000;
   assign mem[5359] = 32'b11111100010111101000010000000100;
   assign mem[5360] = 32'b00000101010101011011110100000000;
   assign mem[5361] = 32'b11111101011011100100001101111100;
   assign mem[5362] = 32'b00000110111011011101001101001000;
   assign mem[5363] = 32'b11111101111101100011100001110000;
   assign mem[5364] = 32'b00000001101111011111110000101100;
   assign mem[5365] = 32'b11110101000100111011111010110000;
   assign mem[5366] = 32'b11101100000110011000110001100000;
   assign mem[5367] = 32'b00000000011101000001000110010001;
   assign mem[5368] = 32'b00000100001001111010000010000000;
   assign mem[5369] = 32'b11111101011101111001111111001100;
   assign mem[5370] = 32'b11111001011111100111110111011000;
   assign mem[5371] = 32'b00000100000010000111111010100000;
   assign mem[5372] = 32'b11111111101010101100111000010100;
   assign mem[5373] = 32'b00000100110010001111001100111000;
   assign mem[5374] = 32'b00000001111100101011010000010100;
   assign mem[5375] = 32'b11110100101110101100100011000000;
   assign mem[5376] = 32'b11111111011100110011011101101100;
   assign mem[5377] = 32'b00000010110011000011011111010000;
   assign mem[5378] = 32'b11111001111001000010101010110000;
   assign mem[5379] = 32'b11111101100110011100101111011000;
   assign mem[5380] = 32'b11111110111010111010111001110000;
   assign mem[5381] = 32'b00000001001111011110100000000110;
   assign mem[5382] = 32'b00000010100111010101000101000100;
   assign mem[5383] = 32'b11111101010001110011010000110000;
   assign mem[5384] = 32'b00000011100101111111101111111000;
   assign mem[5385] = 32'b11110010000011101011001000100000;
   assign mem[5386] = 32'b11111100010101110110101000010100;
   assign mem[5387] = 32'b00000101110100010000100101111000;
   assign mem[5388] = 32'b00000011100010110001010011100100;
   assign mem[5389] = 32'b11111110001011111101000010111010;
   assign mem[5390] = 32'b11110001100100010111100110100000;
   assign mem[5391] = 32'b00010001111000100110011001100000;
   assign mem[5392] = 32'b11111010101010000100101110110000;
   assign mem[5393] = 32'b11110101011101110101100111100000;
   assign mem[5394] = 32'b00000101011011100011101101111000;
   assign mem[5395] = 32'b00001010001010101011111110010000;
   assign mem[5396] = 32'b00001010010101000000011101110000;
   assign mem[5397] = 32'b11111111101001010010111000100011;
   assign mem[5398] = 32'b11111010010001100110111101101000;
   assign mem[5399] = 32'b11110110001001000000010101000000;
   assign mem[5400] = 32'b11111000111000111000110011111000;
   assign mem[5401] = 32'b11101011000110100010011111000000;
   assign mem[5402] = 32'b11111010001100110100110011001000;
   assign mem[5403] = 32'b00000110010011100110110110010000;
   assign mem[5404] = 32'b11110111011010110100101100100000;
   assign mem[5405] = 32'b00000111110001110001011110011000;
   assign mem[5406] = 32'b11111110110101101000100011011010;
   assign mem[5407] = 32'b00000000101101100101100110011011;
   assign mem[5408] = 32'b00001001010111110000101011100000;
   assign mem[5409] = 32'b00000101110110110000001110111000;
   assign mem[5410] = 32'b00000000101110000111000100111100;
   assign mem[5411] = 32'b11111011011010100000110110100000;
   assign mem[5412] = 32'b11111101100101001000011110001100;
   assign mem[5413] = 32'b00000001001101001110011101010110;
   assign mem[5414] = 32'b11110110111010001110010110000000;
   assign mem[5415] = 32'b11111110101100100100011111010100;
   assign mem[5416] = 32'b00000110001001101010110111101000;
   assign mem[5417] = 32'b00000001010001011111101101010010;
   assign mem[5418] = 32'b11111110111010001101000111110110;
   assign mem[5419] = 32'b11111111111011101011101111001010;
   assign mem[5420] = 32'b00000001010101011110110000110000;
   assign mem[5421] = 32'b00000101100101100100011111011000;
   assign mem[5422] = 32'b00000101100101101110011000101000;
   assign mem[5423] = 32'b00000000001001010000011001110011;
   assign mem[5424] = 32'b00000011100110010000011000101100;
   assign mem[5425] = 32'b11110101101010100010001100110000;
   assign mem[5426] = 32'b11111001001101010111001111101000;
   assign mem[5427] = 32'b00000011011101100010000111101000;
   assign mem[5428] = 32'b11111010111010100111101011000000;
   assign mem[5429] = 32'b11111010111001111010001010000000;
   assign mem[5430] = 32'b11111111111001000111101111010100;
   assign mem[5431] = 32'b11110101010110010101100100000000;
   assign mem[5432] = 32'b11111110110100011111011001110100;
   assign mem[5433] = 32'b11111011111111101001100100001000;
   assign mem[5434] = 32'b11101110001001001111111101100000;
   assign mem[5435] = 32'b00001001000110100101110110000000;
   assign mem[5436] = 32'b00000000011011000010101000001111;
   assign mem[5437] = 32'b00000100000010111111000001101000;
   assign mem[5438] = 32'b11111111100010110101101100101001;
   assign mem[5439] = 32'b11111110000111011001001000111100;
   assign mem[5440] = 32'b11111101001001010010010111100100;
   assign mem[5441] = 32'b00000100000010100100100110001000;
   assign mem[5442] = 32'b11110101110000100001011100010000;
   assign mem[5443] = 32'b00000000000100111110011110001110;
   assign mem[5444] = 32'b00000010011111001001011101001000;
   assign mem[5445] = 32'b11111100101001011111110011100000;
   assign mem[5446] = 32'b11111101100011100011110111011100;
   assign mem[5447] = 32'b00000010100100001101000001110100;
   assign mem[5448] = 32'b00000001000000111000100101011010;
   assign mem[5449] = 32'b00000101000100101111100000011000;
   assign mem[5450] = 32'b11111001000000010110010000000000;
   assign mem[5451] = 32'b00000110111101110101001111001000;
   assign mem[5452] = 32'b00000011101000110111101110010100;
   assign mem[5453] = 32'b11110010111111100000111111000000;
   assign mem[5454] = 32'b00000011100000111001011111111100;
   assign mem[5455] = 32'b11111000111011011111000110110000;
   assign mem[5456] = 32'b00000001101101011111111011011010;
   assign mem[5457] = 32'b11111101011101000111100111011000;
   assign mem[5458] = 32'b11111110010110110100100100000000;
   assign mem[5459] = 32'b00000001010110110001000011101000;
   assign mem[5460] = 32'b11111100101011010100110000111000;
   assign mem[5461] = 32'b11110111001000011001011001100000;
   assign mem[5462] = 32'b11111110001011000101111001100010;
   assign mem[5463] = 32'b11111110001011010110011010110100;
   assign mem[5464] = 32'b11110011000000101000111011110000;
   assign mem[5465] = 32'b00000111101010000111001000100000;
   assign mem[5466] = 32'b11111010001111110010101011111000;
   assign mem[5467] = 32'b00000010011100111010111000010000;
   assign mem[5468] = 32'b00000011011000100111001111010000;
   assign mem[5469] = 32'b11111111111111101011001010101110;
   assign mem[5470] = 32'b11110100101001000111111001010000;
   assign mem[5471] = 32'b00000100110100111011001011111000;
   assign mem[5472] = 32'b00000010000100001110000010111100;
   assign mem[5473] = 32'b00000111001010001111100010011000;
   assign mem[5474] = 32'b00000110110011100101011000111000;
   assign mem[5475] = 32'b11111100011111011111111111011000;
   assign mem[5476] = 32'b00000101010111101000100110100000;
   assign mem[5477] = 32'b11111100110101000111000000001100;
   assign mem[5478] = 32'b11111001111011010010101010100000;
   assign mem[5479] = 32'b11110111000011010111010100010000;
   assign mem[5480] = 32'b00000000010101111000100011011101;
   assign mem[5481] = 32'b11111101111110101001111010101100;
   assign mem[5482] = 32'b00000001010111001010011110010100;
   assign mem[5483] = 32'b00000011110100011100101101010100;
   assign mem[5484] = 32'b11110100110010100111011001010000;
   assign mem[5485] = 32'b00000011000001111100011110011100;
   assign mem[5486] = 32'b00000101011000111100010000001000;
   assign mem[5487] = 32'b00000011100001110001100110100000;
   assign mem[5488] = 32'b11111110001000011110001110101000;
   assign mem[5489] = 32'b00000001111000011100101101010110;
   assign mem[5490] = 32'b00000000011101001000110010100000;
   assign mem[5491] = 32'b00000010010111000110110011010100;
   assign mem[5492] = 32'b00000000111110001001101011010010;
   assign mem[5493] = 32'b00000001001000010110001000000000;
   assign mem[5494] = 32'b11111111000110111101110111100100;
   assign mem[5495] = 32'b11111111111111101101001111010001;
   assign mem[5496] = 32'b11111110111011100111011000001110;
   assign mem[5497] = 32'b00000010111100000011001110011100;
   assign mem[5498] = 32'b00000000010000000100101110011001;
   assign mem[5499] = 32'b00000010110100111000001000110100;
   assign mem[5500] = 32'b11111110010011001010110101101010;
   assign mem[5501] = 32'b00001000111010111011100011100000;
   assign mem[5502] = 32'b11111011110001110100111001100000;
   assign mem[5503] = 32'b00000000101000000100101100000000;
   assign mem[5504] = 32'b00000111111000101011011001001000;
   assign mem[5505] = 32'b00000101101100111000000100100000;
   assign mem[5506] = 32'b11110110100000000001010001010000;
   assign mem[5507] = 32'b11111111101101000010100000110101;
   assign mem[5508] = 32'b00000010100111001001000000101100;
   assign mem[5509] = 32'b11111011110000000010001010001000;
   assign mem[5510] = 32'b11110000011001001100100010110000;
   assign mem[5511] = 32'b00001000000000001000100010010000;
   assign mem[5512] = 32'b00000010000111110001101000010100;
   assign mem[5513] = 32'b00000010100101100010000111111000;
   assign mem[5514] = 32'b11110001100010000101100010100000;
   assign mem[5515] = 32'b00000101100011101100011100000000;
   assign mem[5516] = 32'b00000011011010000101000010001000;
   assign mem[5517] = 32'b00000001001001011110001010110110;
   assign mem[5518] = 32'b11111010101001000010110011000000;
   assign mem[5519] = 32'b11111100101011111000010011001000;
   assign mem[5520] = 32'b00000110110011001110011110001000;
   assign mem[5521] = 32'b11111011101011101101110001111000;
   assign mem[5522] = 32'b11111101101101011101000011100000;
   assign mem[5523] = 32'b11111100110000000101000000111100;
   assign mem[5524] = 32'b00000111101101010110110001100000;
   assign mem[5525] = 32'b00000010000000010110111011111100;
   assign mem[5526] = 32'b11111110110111111011101111111000;
   assign mem[5527] = 32'b00000100100111101011001000101000;
   assign mem[5528] = 32'b11111011000101010011101100000000;
   assign mem[5529] = 32'b11111110001011011101110011100100;
   assign mem[5530] = 32'b11111000101101110011000110111000;
   assign mem[5531] = 32'b00000100111010011100011100011000;
   assign mem[5532] = 32'b11111001001111000000001111001000;
   assign mem[5533] = 32'b11111000001001111001000100001000;
   assign mem[5534] = 32'b11111111101100100101100010010000;
   assign mem[5535] = 32'b00001000111011000000000011010000;
   assign mem[5536] = 32'b00000001100101100010011001011010;
   assign mem[5537] = 32'b00000111011001111011110010000000;
   assign mem[5538] = 32'b00000010111101110110010100101100;
   assign mem[5539] = 32'b00000000100000111010111110000111;
   assign mem[5540] = 32'b11111110011000001110001011011100;
   assign mem[5541] = 32'b11110101001001010111001000000000;
   assign mem[5542] = 32'b00000111010011110000001000100000;
   assign mem[5543] = 32'b11110110011010101111100100100000;
   assign mem[5544] = 32'b11110000010000110100111100000000;
   assign mem[5545] = 32'b00000110101100010010101010100000;
   assign mem[5546] = 32'b00001100000111010111110101000000;
   assign mem[5547] = 32'b00000001100010000101100110101110;
   assign mem[5548] = 32'b11110000111011011010100001010000;
   assign mem[5549] = 32'b00000010010001000011001111101100;
   assign mem[5550] = 32'b00000011001110011001101100101000;
   assign mem[5551] = 32'b11111111011001011001001100110110;
   assign mem[5552] = 32'b00000110101101011011000101110000;
   assign mem[5553] = 32'b11111111111011110110010100100001;
   assign mem[5554] = 32'b00000010000111000101010101010000;
   assign mem[5555] = 32'b11101100011010101001101100100000;
   assign mem[5556] = 32'b11110101111000100110110100110000;
   assign mem[5557] = 32'b11111101110110010010000100101100;
   assign mem[5558] = 32'b00000000010100001111011011100111;
   assign mem[5559] = 32'b11111110101100000110001001100100;
   assign mem[5560] = 32'b11111000010111001010110100100000;
   assign mem[5561] = 32'b00001010101010110000111010100000;
   assign mem[5562] = 32'b11111010100110010100011001100000;
   assign mem[5563] = 32'b00001011110111110011011010000000;
   assign mem[5564] = 32'b00000101001110001011001001001000;
   assign mem[5565] = 32'b00000001011110111111101000001000;
   assign mem[5566] = 32'b11101110111011101011100111100000;
   assign mem[5567] = 32'b11101111100011001101011010000000;
   assign mem[5568] = 32'b11111101111010000101111100100000;
   assign mem[5569] = 32'b00000100100001000111010010010000;
   assign mem[5570] = 32'b00000010001110011011000100011000;
   assign mem[5571] = 32'b11111100100001110111100000101000;
   assign mem[5572] = 32'b00000100111000110001011000001000;
   assign mem[5573] = 32'b00000001010101101010001101110000;
   assign mem[5574] = 32'b11111100000010111011010011111100;
   assign mem[5575] = 32'b11110110000101100111001110110000;
   assign mem[5576] = 32'b11111100011010000100110000000100;
   assign mem[5577] = 32'b00000011011001111011111111000000;
   assign mem[5578] = 32'b00000100101010001100011111101000;
   assign mem[5579] = 32'b00000001111100000111000001010110;
   assign mem[5580] = 32'b11111011101100101011111111000000;
   assign mem[5581] = 32'b11111100100100001001010111111000;
   assign mem[5582] = 32'b00000010000101101001001011101100;
   assign mem[5583] = 32'b00000010001001010000000111111000;
   assign mem[5584] = 32'b00000001000001001110100101101110;
   assign mem[5585] = 32'b11111001011111110101000010100000;
   assign mem[5586] = 32'b11111010111100010011010011111000;
   assign mem[5587] = 32'b00000101010101101000010010011000;
   assign mem[5588] = 32'b11111101101011101110101111000000;
   assign mem[5589] = 32'b00000000010100010001110100010001;
   assign mem[5590] = 32'b00000010010011010000101111011000;
   assign mem[5591] = 32'b11111110111010010001111111010010;
   assign mem[5592] = 32'b00000011101110010101111111100100;
   assign mem[5593] = 32'b11111101000011100110101000101100;
   assign mem[5594] = 32'b00000011001100001000100110110100;
   assign mem[5595] = 32'b11111111101111101100011101011101;
   assign mem[5596] = 32'b00000000101100110101001001110010;
   assign mem[5597] = 32'b11111111011000111110101011000110;
   assign mem[5598] = 32'b00000001111000001001010000010110;
   assign mem[5599] = 32'b00000000000011010011001111100110;
   assign mem[5600] = 32'b00000010000001111010100100001000;
   assign mem[5601] = 32'b00000101111000110000110001010000;
   assign mem[5602] = 32'b11110110011011000000101001000000;
   assign mem[5603] = 32'b00000011100011100010110110110100;
   assign mem[5604] = 32'b11110110011001011110010100000000;
   assign mem[5605] = 32'b00000101000101000101001010101000;
   assign mem[5606] = 32'b11111101001101101101100110111100;
   assign mem[5607] = 32'b00000001010101011010011000100110;
   assign mem[5608] = 32'b11111100001101010100011010001000;
   assign mem[5609] = 32'b11111110111100010000100000001100;
   assign mem[5610] = 32'b11110110111010100010001110110000;
   assign mem[5611] = 32'b00001010010101111101000110000000;
   assign mem[5612] = 32'b11111000001000011001111001101000;
   assign mem[5613] = 32'b11110001111111001011011100100000;
   assign mem[5614] = 32'b00001000001000010101100001000000;
   assign mem[5615] = 32'b00000100111101100010011011110000;
   assign mem[5616] = 32'b00001111010011010101100011000000;
   assign mem[5617] = 32'b00000100010010010100101001100000;
   assign mem[5618] = 32'b11111000100111010100011111110000;
   assign mem[5619] = 32'b11111011010101101001010110101000;
   assign mem[5620] = 32'b11111010111101001110011011011000;
   assign mem[5621] = 32'b11110100110011010110101100100000;
   assign mem[5622] = 32'b00000001011010011100100011111110;
   assign mem[5623] = 32'b00000111101001100110101111001000;
   assign mem[5624] = 32'b11111110111101111011001000010000;
   assign mem[5625] = 32'b11110100110100001000101100110000;
   assign mem[5626] = 32'b11111101100011011001110000110000;
   assign mem[5627] = 32'b00000110110111001101111101011000;
   assign mem[5628] = 32'b00000110000101101101100011011000;
   assign mem[5629] = 32'b00000111001111111000001000010000;
   assign mem[5630] = 32'b00000110110101100010101110111000;
   assign mem[5631] = 32'b00001100011110100101110100100000;
   assign mem[5632] = 32'b00001001001010111001010010010000;
   assign mem[5633] = 32'b11110000010010011100011110000000;
   assign mem[5634] = 32'b11111111001111010111100111100111;
   assign mem[5635] = 32'b11101000100011000110011010000000;
   assign mem[5636] = 32'b11111010111101110111110000010000;
   assign mem[5637] = 32'b00000000110011111100000100110010;
   assign mem[5638] = 32'b11111110010010000010010001100010;
   assign mem[5639] = 32'b11111111011011000100000101001010;
   assign mem[5640] = 32'b00000001000110100000110010010110;
   assign mem[5641] = 32'b11110101010001000001110111000000;
   assign mem[5642] = 32'b11111100111011001100001010100100;
   assign mem[5643] = 32'b00000010001111110001000000100000;
   assign mem[5644] = 32'b11111100100001111111010101111100;
   assign mem[5645] = 32'b00001000101000100010000010100000;
   assign mem[5646] = 32'b11110111111111100000010101100000;
   assign mem[5647] = 32'b00000100000101110010010000001000;
   assign mem[5648] = 32'b11111110010010000110111110010110;
   assign mem[5649] = 32'b00000001101011101011010001011100;
   assign mem[5650] = 32'b11111101011011000100011010100000;
   assign mem[5651] = 32'b11110110110001111100110000000000;
   assign mem[5652] = 32'b11111100100101001100010111111000;
   assign mem[5653] = 32'b00001000100100001011000011010000;
   assign mem[5654] = 32'b11110010010010111100101010110000;
   assign mem[5655] = 32'b00001001000101011000000001110000;
   assign mem[5656] = 32'b11111100111101001110000110011100;
   assign mem[5657] = 32'b00000101010011011101010111001000;
   assign mem[5658] = 32'b00000011001110101111001010001000;
   assign mem[5659] = 32'b11111101010101111111000000011100;
   assign mem[5660] = 32'b11111101000001111001000001100100;
   assign mem[5661] = 32'b00000000001111100101001011001101;
   assign mem[5662] = 32'b11111010100000011011111111101000;
   assign mem[5663] = 32'b11111111110100000110001010010100;
   assign mem[5664] = 32'b11111010010101111110101001100000;
   assign mem[5665] = 32'b00000110110101100100100001100000;
   assign mem[5666] = 32'b00000100111000100010101001011000;
   assign mem[5667] = 32'b00000110111110100000110101110000;
   assign mem[5668] = 32'b11111001011110101110001111011000;
   assign mem[5669] = 32'b11111001000001111110101011100000;
   assign mem[5670] = 32'b00000110111010101110101111100000;
   assign mem[5671] = 32'b11111101110011110110100110010000;
   assign mem[5672] = 32'b00000001100111010101100010010100;
   assign mem[5673] = 32'b00000000010010011100011000100110;
   assign mem[5674] = 32'b00000111101101010001001000101000;
   assign mem[5675] = 32'b11110000110110011000011111110000;
   assign mem[5676] = 32'b00000011111010011010000011001000;
   assign mem[5677] = 32'b00000001000010000011101111011010;
   assign mem[5678] = 32'b11111100011000010000010001100000;
   assign mem[5679] = 32'b11111100101111000101011100110100;
   assign mem[5680] = 32'b00000101000000100000001111111000;
   assign mem[5681] = 32'b00000110011001001100110000001000;
   assign mem[5682] = 32'b00000110011101101111100110010000;
   assign mem[5683] = 32'b00000111001100000111101100100000;
   assign mem[5684] = 32'b11111011101110001100011111000000;
   assign mem[5685] = 32'b11101111010111110010100011100000;
   assign mem[5686] = 32'b11110110100000100110111110110000;
   assign mem[5687] = 32'b00000010101000101000011000001100;
   assign mem[5688] = 32'b11111101011111100001111011011100;
   assign mem[5689] = 32'b00000110111110010101000110100000;
   assign mem[5690] = 32'b11111110111010101110110001100000;
   assign mem[5691] = 32'b11110000001010110010000111100000;
   assign mem[5692] = 32'b00000100010111101101001010011000;
   assign mem[5693] = 32'b00000001011101011010001111100100;
   assign mem[5694] = 32'b11111000110101010001111011110000;
   assign mem[5695] = 32'b11111101111100001011000110010000;
   assign mem[5696] = 32'b11111110010001101100011001001000;
   assign mem[5697] = 32'b00000100100111110001010111110000;
   assign mem[5698] = 32'b11111110101101110001000101010110;
   assign mem[5699] = 32'b00000000001000001000101111111000;
   assign mem[5700] = 32'b00000110101010000010011001011000;
   assign mem[5701] = 32'b11111110100110000101111100100000;
   assign mem[5702] = 32'b00001001100001000001110000000000;
   assign mem[5703] = 32'b11111110001110001010011110110000;
   assign mem[5704] = 32'b11111101110100101110100011100000;
   assign mem[5705] = 32'b11111100000101111010001001101000;
   assign mem[5706] = 32'b11111101110000000101011101010100;
   assign mem[5707] = 32'b00000001000111101101000010101100;
   assign mem[5708] = 32'b11111000011000101010001010010000;
   assign mem[5709] = 32'b00000010010010101000100111111000;
   assign mem[5710] = 32'b00000111011100111001100000000000;
   assign mem[5711] = 32'b11111101010010010100010111011100;
   assign mem[5712] = 32'b00000001010000100111011001111010;
   assign mem[5713] = 32'b00000010101110100101010000100100;
   assign mem[5714] = 32'b11111111010001010000000101100001;
   assign mem[5715] = 32'b11111010011101000101000110111000;
   assign mem[5716] = 32'b11110101000110100100100010100000;
   assign mem[5717] = 32'b11111111101011010100111000010001;
   assign mem[5718] = 32'b00000010110101111111111011010000;
   assign mem[5719] = 32'b00000100011111010010110110100000;
   assign mem[5720] = 32'b11111101101101000010110001000000;
   assign mem[5721] = 32'b00010000011100010110000111000000;
   assign mem[5722] = 32'b11110111001000110010010110010000;
   assign mem[5723] = 32'b11110101101010111101101001010000;
   assign mem[5724] = 32'b11111110100010110000111000100010;
   assign mem[5725] = 32'b00000110011110100000111010000000;
   assign mem[5726] = 32'b00001010000100001000001011100000;
   assign mem[5727] = 32'b00000110000001100100001110000000;
   assign mem[5728] = 32'b11111000010101100000111100011000;
   assign mem[5729] = 32'b11111100110100010001101101110000;
   assign mem[5730] = 32'b11111110100101011111100101011110;
   assign mem[5731] = 32'b00010000011101001111011011000000;
   assign mem[5732] = 32'b11110111101010100110100010000000;
   assign mem[5733] = 32'b11110001010010110101111111100000;
   assign mem[5734] = 32'b00000111101101110110011111011000;
   assign mem[5735] = 32'b00000011110100100101001011110000;
   assign mem[5736] = 32'b00001001110101101000011101100000;
   assign mem[5737] = 32'b11111111100011101010110110101100;
   assign mem[5738] = 32'b11111001100000011100011111010000;
   assign mem[5739] = 32'b11111001111101010110010111101000;
   assign mem[5740] = 32'b00000000010001001110011010111101;
   assign mem[5741] = 32'b00001100111100011101100100010000;
   assign mem[5742] = 32'b00000110001111110001110111010000;
   assign mem[5743] = 32'b11100101001010001000110000100000;
   assign mem[5744] = 32'b00001101000000010100010001110000;
   assign mem[5745] = 32'b11101110000010111111101110100000;
   assign mem[5746] = 32'b11111111001001110101110110000100;
   assign mem[5747] = 32'b11110010110011001100101001000000;
   assign mem[5748] = 32'b11110111010110010101100110000000;
   assign mem[5749] = 32'b11110111110011010110100101000000;
   assign mem[5750] = 32'b11111001101011110110010101100000;
   assign mem[5751] = 32'b00001001101100001011110101110000;
   assign mem[5752] = 32'b11111111001000011101110110010110;
   assign mem[5753] = 32'b00000001011110100001010010111100;
   assign mem[5754] = 32'b00001001110100100010110000000000;
   assign mem[5755] = 32'b11101111001011011011100111100000;
   assign mem[5756] = 32'b11111100000111000101100110111000;
   assign mem[5757] = 32'b11111111000100100111000010000101;
   assign mem[5758] = 32'b00000100100011010010000001111000;
   assign mem[5759] = 32'b11111110111111010101011100000010;
   assign mem[5760] = 32'b11111101010001000010100000110100;
   assign mem[5761] = 32'b11111101001111010100111111111000;
   assign mem[5762] = 32'b11111101001001101110111101100100;
   assign mem[5763] = 32'b00000010011110010010110110001000;
   assign mem[5764] = 32'b00001111011111000100011110110000;
   assign mem[5765] = 32'b11111111100011100010111001001101;
   assign mem[5766] = 32'b00001010101110000100001100110000;
   assign mem[5767] = 32'b11110100010110000111110100010000;
   assign mem[5768] = 32'b00000000110101000100100010110011;
   assign mem[5769] = 32'b11101111100001111110001101000000;
   assign mem[5770] = 32'b00000011010000001110111000000000;
   assign mem[5771] = 32'b11111011000111110100001101010000;
   assign mem[5772] = 32'b11111111011101000101011010000111;
   assign mem[5773] = 32'b11111111100011010001010100000001;
   assign mem[5774] = 32'b00000001010101110110001101100110;
   assign mem[5775] = 32'b11110101010010010110000110110000;
   assign mem[5776] = 32'b11111101100111001111010000101000;
   assign mem[5777] = 32'b00000000100100100101010011110111;
   assign mem[5778] = 32'b00000001010011111101100001000110;
   assign mem[5779] = 32'b11111111111100101100100011011011;
   assign mem[5780] = 32'b00001000100010100010011100110000;
   assign mem[5781] = 32'b11111010010100010111010110010000;
   assign mem[5782] = 32'b11111100100010110010110010101000;
   assign mem[5783] = 32'b11111100110101100011110000000000;
   assign mem[5784] = 32'b11110010011110010101111001100000;
   assign mem[5785] = 32'b11111100001010111001000001010000;
   assign mem[5786] = 32'b00000001100001101100110001100110;
   assign mem[5787] = 32'b11111110001000111111110100011010;
   assign mem[5788] = 32'b00001001011011001011100011000000;
   assign mem[5789] = 32'b00000100100001001000111110000000;
   assign mem[5790] = 32'b00000100000010010010100000101000;
   assign mem[5791] = 32'b11110010000000100000110001000000;
   assign mem[5792] = 32'b11110101101111110111111000000000;
   assign mem[5793] = 32'b11110010011100001100101011100000;
   assign mem[5794] = 32'b11110000000101010011100101010000;
   assign mem[5795] = 32'b00001110001010011110110110000000;
   assign mem[5796] = 32'b00000010100101101000110011110100;
   assign mem[5797] = 32'b11101101101101111111110011100000;
   assign mem[5798] = 32'b00000100011110010001101000001000;
   assign mem[5799] = 32'b00000110011100101110100010000000;
   assign mem[5800] = 32'b11110010000100101000111010010000;
   assign mem[5801] = 32'b11111010101011101100110100111000;
   assign mem[5802] = 32'b11101001000100001110100001000000;
   assign mem[5803] = 32'b11110001001111010110010101110000;
   assign mem[5804] = 32'b11111100000110110110101110100000;
   assign mem[5805] = 32'b00001100000111010101110010100000;
   assign mem[5806] = 32'b00010001000001011011110111000000;
   assign mem[5807] = 32'b11111101100010001111000101000000;
   assign mem[5808] = 32'b00000000000100110000110111011010;
   assign mem[5809] = 32'b11110111000000110001101100000000;
   assign mem[5810] = 32'b11111101101101000011110111111100;
   assign mem[5811] = 32'b00000110001100101001011100000000;
   assign mem[5812] = 32'b00000000011001101110000010100101;
   assign mem[5813] = 32'b00000111001100000101110001110000;
   assign mem[5814] = 32'b00001001000000111011101001000000;
   assign mem[5815] = 32'b11110010001011001110100001100000;
   assign mem[5816] = 32'b00000001000001001010010110110010;
   assign mem[5817] = 32'b11111000110101000001101011001000;
   assign mem[5818] = 32'b00000010000100011011000010100100;
   assign mem[5819] = 32'b11111011100100100000110001110000;
   assign mem[5820] = 32'b11110101101101000110110101000000;
   assign mem[5821] = 32'b11111111110001010110000011000110;
   assign mem[5822] = 32'b11111011100111010000001001111000;
   assign mem[5823] = 32'b00000100001000111011101010110000;
   assign mem[5824] = 32'b00000000001000011000101100110101;
   assign mem[5825] = 32'b11111101000110110101000101100000;
   assign mem[5826] = 32'b11111111101010011111111000001110;
   assign mem[5827] = 32'b11111111100010101100000110111111;
   assign mem[5828] = 32'b00000000101000001000010110101111;
   assign mem[5829] = 32'b00000000110000101101100110101010;
   assign mem[5830] = 32'b11110010001111001000010101010000;
   assign mem[5831] = 32'b11111111110100101010100101011011;
   assign mem[5832] = 32'b11111111010011100010100101010001;
   assign mem[5833] = 32'b00000010101100100101011011100000;
   assign mem[5834] = 32'b00000110001011011101101101010000;
   assign mem[5835] = 32'b00000010001000111001010000010100;
   assign mem[5836] = 32'b11111101101100000010000111011100;
   assign mem[5837] = 32'b00000111101100000111111010000000;
   assign mem[5838] = 32'b00000000110101000001000100000111;
   assign mem[5839] = 32'b11110111101000011000000000100000;
   assign mem[5840] = 32'b00000000010110001010001101001001;
   assign mem[5841] = 32'b11111010110101101010101010100000;
   assign mem[5842] = 32'b11111110000000110100001110000110;
   assign mem[5843] = 32'b11111100101110100011010011101000;
   assign mem[5844] = 32'b11111100101110011111100111110100;
   assign mem[5845] = 32'b00000000000111110100101101011111;
   assign mem[5846] = 32'b00001011000100110001100010100000;
   assign mem[5847] = 32'b00000011111111010001100111011000;
   assign mem[5848] = 32'b11111011001011011001010100111000;
   assign mem[5849] = 32'b11111010101100101111000111101000;
   assign mem[5850] = 32'b11111110111010100001000001110000;
   assign mem[5851] = 32'b00001001010011100100001001100000;
   assign mem[5852] = 32'b11111110111110011111001111010010;
   assign mem[5853] = 32'b00000000001111011110111000100100;
   assign mem[5854] = 32'b00000001011000100011000101110000;
   assign mem[5855] = 32'b00000000011101000101001101001010;
   assign mem[5856] = 32'b11111011001001110111110001011000;
   assign mem[5857] = 32'b00000011000111010110000001110000;
   assign mem[5858] = 32'b11111000000010010010110100010000;
   assign mem[5859] = 32'b11101100100011011001000101000000;
   assign mem[5860] = 32'b11111000110011001101110100010000;
   assign mem[5861] = 32'b11110010101100100100000111010000;
   assign mem[5862] = 32'b11101101010110111111000111100000;
   assign mem[5863] = 32'b11110011001111000001001010010000;
   assign mem[5864] = 32'b00000001010100100110101011000010;
   assign mem[5865] = 32'b00001010101111011010100011010000;
   assign mem[5866] = 32'b11111011101101000110001111110000;
   assign mem[5867] = 32'b00000000101011000101101010100001;
   assign mem[5868] = 32'b00000100001010110011101101101000;
   assign mem[5869] = 32'b11111101100111000000010111011000;
   assign mem[5870] = 32'b00001001111001100110011110110000;
   assign mem[5871] = 32'b11110111101110110100000011100000;
   assign mem[5872] = 32'b11111101000001111110001010110100;
   assign mem[5873] = 32'b11110000110100011001111101010000;
   assign mem[5874] = 32'b11111001011000100001001101100000;
   assign mem[5875] = 32'b11111111011111111010110001001001;
   assign mem[5876] = 32'b00000011111011110001010111111000;
   assign mem[5877] = 32'b11111101111101000111010001110000;
   assign mem[5878] = 32'b00000111010101111010100110101000;
   assign mem[5879] = 32'b00000011111011000010010010111000;
   assign mem[5880] = 32'b11111010001110011110101001110000;
   assign mem[5881] = 32'b11110110111101011001001111100000;
   assign mem[5882] = 32'b00000001010001000110000100000100;
   assign mem[5883] = 32'b00000111011011001111011010111000;
   assign mem[5884] = 32'b00000111100000011000000110110000;
   assign mem[5885] = 32'b00000110001000010000011110010000;
   assign mem[5886] = 32'b00000101100110111101001010011000;
   assign mem[5887] = 32'b00000000111011011101011001011010;
   assign mem[5888] = 32'b11111101010000010100010011011000;
   assign mem[5889] = 32'b11101101000110000111000110000000;
   assign mem[5890] = 32'b00000010100001101010110101101000;
   assign mem[5891] = 32'b11110101100010001111010000100000;
   assign mem[5892] = 32'b11111100000001011000011111000000;
   assign mem[5893] = 32'b11111110001110001010100001011100;
   assign mem[5894] = 32'b11111001010111011001011011100000;
   assign mem[5895] = 32'b11111011111000011100001000100000;
   assign mem[5896] = 32'b00001010100011010001000000000000;
   assign mem[5897] = 32'b00000000001011010011101010000010;
   assign mem[5898] = 32'b00000010111001110011010110110000;
   assign mem[5899] = 32'b11111111001010101000100111011100;
   assign mem[5900] = 32'b00000000000001100001101100110111;
   assign mem[5901] = 32'b00000110000101010011011111001000;
   assign mem[5902] = 32'b11111011101010101011100000100000;
   assign mem[5903] = 32'b00001000110011010001110101100000;
   assign mem[5904] = 32'b00000101101111011011111011001000;
   assign mem[5905] = 32'b00000111111111010111011001000000;
   assign mem[5906] = 32'b11111101100110101101011011010000;
   assign mem[5907] = 32'b11111101111111000100011110011100;
   assign mem[5908] = 32'b11111011000010110001101000001000;
   assign mem[5909] = 32'b11111011110111111100110110100000;
   assign mem[5910] = 32'b00000101011110011000010000100000;
   assign mem[5911] = 32'b11111100010111111010101100001100;
   assign mem[5912] = 32'b00001001100000001011001110010000;
   assign mem[5913] = 32'b11111100110000100010100100111100;
   assign mem[5914] = 32'b00001000110001110111010011110000;
   assign mem[5915] = 32'b11101010011001111001011100100000;
   assign mem[5916] = 32'b11110100010010011011001001110000;
   assign mem[5917] = 32'b11111000000010011100010001010000;
   assign mem[5918] = 32'b00001000100001111110100010100000;
   assign mem[5919] = 32'b11110100110100010110001101010000;
   assign mem[5920] = 32'b11110110000110011111110011000000;
   assign mem[5921] = 32'b11111100000010100011111010001100;
   assign mem[5922] = 32'b11110011111100110010001001110000;
   assign mem[5923] = 32'b11111010010010100100111111011000;
   assign mem[5924] = 32'b00000010101010011100100000001100;
   assign mem[5925] = 32'b00001110000011101110010101010000;
   assign mem[5926] = 32'b00000000101110101110111110100001;
   assign mem[5927] = 32'b00001100001111101111001101100000;
   assign mem[5928] = 32'b11111111110010000100011010100111;
   assign mem[5929] = 32'b11111100010100001111101100111000;
   assign mem[5930] = 32'b00000100100001011100111011001000;
   assign mem[5931] = 32'b11111100001010000010100011011100;
   assign mem[5932] = 32'b11111010111000011101011100011000;
   assign mem[5933] = 32'b11111011000011101001011010000000;
   assign mem[5934] = 32'b11110101000111100010100001000000;
   assign mem[5935] = 32'b00000100111100010010110000100000;
   assign mem[5936] = 32'b11111110100011001010000110011000;
   assign mem[5937] = 32'b00000101110000100111101100000000;
   assign mem[5938] = 32'b00000100110111010110001110111000;
   assign mem[5939] = 32'b11111110110111010011010111111110;
   assign mem[5940] = 32'b11111011111000111011010111010000;
   assign mem[5941] = 32'b11110100110010010010110010100000;
   assign mem[5942] = 32'b11111010111101111111011000101000;
   assign mem[5943] = 32'b11111100101101001111101000111000;
   assign mem[5944] = 32'b11111111100010110000110101100100;
   assign mem[5945] = 32'b00001000100011010110010000000000;
   assign mem[5946] = 32'b00000111001111111000111110110000;
   assign mem[5947] = 32'b11111001011000011010111111101000;
   assign mem[5948] = 32'b11111110101001100101011101001010;
   assign mem[5949] = 32'b00000101010011010111110111010000;
   assign mem[5950] = 32'b11111001111001010001001101001000;
   assign mem[5951] = 32'b11101010010111010000000101100000;
   assign mem[5952] = 32'b11111100010001011110000110011100;
   assign mem[5953] = 32'b00000101101011011101001011001000;
   assign mem[5954] = 32'b11111000011101101101100100100000;
   assign mem[5955] = 32'b00000001000011000110111000000000;
   assign mem[5956] = 32'b00001000111100010011000111110000;
   assign mem[5957] = 32'b11111111110011111111001001111001;
   assign mem[5958] = 32'b00000011001001100000100011000100;
   assign mem[5959] = 32'b11111111100101010111001100000101;
   assign mem[5960] = 32'b00000100001100110011011010111000;
   assign mem[5961] = 32'b11111101011110011101111100001100;
   assign mem[5962] = 32'b00000010010110111111100001000100;
   assign mem[5963] = 32'b11111011000110111011010100100000;
   assign mem[5964] = 32'b00001000101101000111010101100000;
   assign mem[5965] = 32'b11110100100110010011101110100000;
   assign mem[5966] = 32'b11110110110101001001011010010000;
   assign mem[5967] = 32'b11110100111111100111100001110000;
   assign mem[5968] = 32'b00000100110000101111100100010000;
   assign mem[5969] = 32'b11111100000111001011110100010000;
   assign mem[5970] = 32'b00000000011100011010000011011100;
   assign mem[5971] = 32'b11110111101001001100001000100000;
   assign mem[5972] = 32'b11111110101101100001110101001010;
   assign mem[5973] = 32'b00000001101000011011100101011000;
   assign mem[5974] = 32'b00000110001000010100111101001000;
   assign mem[5975] = 32'b00000001000111101100100111100100;
   assign mem[5976] = 32'b11111101101101110101110011111100;
   assign mem[5977] = 32'b11111101010100101111101000001000;
   assign mem[5978] = 32'b00000010111111111011001000100000;
   assign mem[5979] = 32'b11111101110100010011101011111000;
   assign mem[5980] = 32'b11110101111000010101100101010000;
   assign mem[5981] = 32'b00000001101110010001011111100110;
   assign mem[5982] = 32'b00000011011101100110010011001000;
   assign mem[5983] = 32'b00000100110110111110010000100000;
   assign mem[5984] = 32'b00000011000101100000111100111100;
   assign mem[5985] = 32'b11101101100101010000010101000000;
   assign mem[5986] = 32'b11110100101000101100101101100000;
   assign mem[5987] = 32'b00000101100110100110100001101000;
   assign mem[5988] = 32'b00000101100100111110110110000000;
   assign mem[5989] = 32'b11111111110110000000101001101111;
   assign mem[5990] = 32'b00000111001101001100100010010000;
   assign mem[5991] = 32'b11111101111100001001111111100000;
   assign mem[5992] = 32'b11111111100010110110101110100000;
   assign mem[5993] = 32'b11111101001001000011010101000000;
   assign mem[5994] = 32'b00000001110010110110111110011000;
   assign mem[5995] = 32'b11110001000011110101110111010000;
   assign mem[5996] = 32'b11110101101110110011011111110000;
   assign mem[5997] = 32'b11111011110001111010101011000000;
   assign mem[5998] = 32'b00000011100100100111000101000000;
   assign mem[5999] = 32'b00000100000001101000010101000000;
   assign mem[6000] = 32'b00001011001101101011001000110000;
   assign mem[6001] = 32'b11111110110100110011101001101010;
   assign mem[6002] = 32'b00000000011001100000001101010110;
   assign mem[6003] = 32'b11110110110001110000100001010000;
   assign mem[6004] = 32'b00000110110110011100101001111000;
   assign mem[6005] = 32'b11101100000011000010101011100000;
   assign mem[6006] = 32'b11111101001100101111101111010100;
   assign mem[6007] = 32'b11111101000010101011110111100000;
   assign mem[6008] = 32'b00000111011110111111011111001000;
   assign mem[6009] = 32'b11111100110100100100101100010000;
   assign mem[6010] = 32'b11111101010101111100011100110000;
   assign mem[6011] = 32'b11111101110111001010111001010100;
   assign mem[6012] = 32'b11111111000011100011010101110101;
   assign mem[6013] = 32'b00000010001001100111010001000100;
   assign mem[6014] = 32'b11111111100001101110011001000000;
   assign mem[6015] = 32'b11111010011001111010000111001000;
   assign mem[6016] = 32'b11111010110011101111110100011000;
   assign mem[6017] = 32'b00000011001000101111110011100100;
   assign mem[6018] = 32'b00000000011100011010010100001101;
   assign mem[6019] = 32'b00000001100010001111111100100100;
   assign mem[6020] = 32'b00000100000011000001101100010000;
   assign mem[6021] = 32'b00000001001011101101110001101000;
   assign mem[6022] = 32'b00000001001010011100111111001100;
   assign mem[6023] = 32'b00000000110111001000100001101000;
   assign mem[6024] = 32'b00000011000110110010000001110000;
   assign mem[6025] = 32'b11110010111111000101010001110000;
   assign mem[6026] = 32'b11101011000111010111010011100000;
   assign mem[6027] = 32'b11111101010101111000110011010100;
   assign mem[6028] = 32'b00000000100100010001100110111100;
   assign mem[6029] = 32'b00000011011000101101101110101000;
   assign mem[6030] = 32'b11100110011111100000011101000000;
   assign mem[6031] = 32'b00001000101001000110100101110000;
   assign mem[6032] = 32'b11110101111010111111110000100000;
   assign mem[6033] = 32'b11111001111000011010000000001000;
   assign mem[6034] = 32'b00000100000011011000001111001000;
   assign mem[6035] = 32'b00001010000111100100011011110000;
   assign mem[6036] = 32'b00000101001110101011001100100000;
   assign mem[6037] = 32'b00001010110001100101011100000000;
   assign mem[6038] = 32'b11111111000001001101101110111000;
   assign mem[6039] = 32'b11101011100011000110000111100000;
   assign mem[6040] = 32'b11110111111001100111110011100000;
   assign mem[6041] = 32'b11111001011111011110001000000000;
   assign mem[6042] = 32'b11111101010010011001110101100000;
   assign mem[6043] = 32'b00000100011111100110010010010000;
   assign mem[6044] = 32'b11111111100101011011101011010100;
   assign mem[6045] = 32'b00000111000000100111100100101000;
   assign mem[6046] = 32'b11110111111010110010001100100000;
   assign mem[6047] = 32'b11111111110100000001010101010110;
   assign mem[6048] = 32'b00000011011110101011000101000000;
   assign mem[6049] = 32'b11111100110101110011111100110100;
   assign mem[6050] = 32'b00000100000110111111010110010000;
   assign mem[6051] = 32'b11110010110101101010100100110000;
   assign mem[6052] = 32'b11111101011001111110010011001000;
   assign mem[6053] = 32'b11111100001100110111110110010100;
   assign mem[6054] = 32'b11110011100100000011100001100000;
   assign mem[6055] = 32'b00000010110001011001001000001100;
   assign mem[6056] = 32'b00001001101011110011100010110000;
   assign mem[6057] = 32'b00000000110101000101000101100110;
   assign mem[6058] = 32'b00000010000000101011100010001000;
   assign mem[6059] = 32'b11111010110001001101111101001000;
   assign mem[6060] = 32'b00000111001011100011001000000000;
   assign mem[6061] = 32'b11110111001101000101011110000000;
   assign mem[6062] = 32'b00000101110010010000000011011000;
   assign mem[6063] = 32'b11111100110001101010000011110100;
   assign mem[6064] = 32'b00000000010101010011100101111111;
   assign mem[6065] = 32'b11110001001110110001111010110000;
   assign mem[6066] = 32'b11101110000001001110100001000000;
   assign mem[6067] = 32'b00000100001110111000011000010000;
   assign mem[6068] = 32'b00000100111111110100001001011000;
   assign mem[6069] = 32'b00000010001110100101111101011000;
   assign mem[6070] = 32'b00000010100010001010011101000000;
   assign mem[6071] = 32'b11111000111001111100100100010000;
   assign mem[6072] = 32'b11101001001101001110010110000000;
   assign mem[6073] = 32'b11111000011101010100111011100000;
   assign mem[6074] = 32'b00000000000010110110100101101001;
   assign mem[6075] = 32'b00001011011000010000110010100000;
   assign mem[6076] = 32'b00000011101101010000010010011100;
   assign mem[6077] = 32'b11111010011100111001001000111000;
   assign mem[6078] = 32'b11111111110101100101010000000000;
   assign mem[6079] = 32'b11111100111100101010100000111100;
   assign mem[6080] = 32'b11111110011000101101110010010110;
   assign mem[6081] = 32'b00000111111110101001110001011000;
   assign mem[6082] = 32'b11110001010001010010000100100000;
   assign mem[6083] = 32'b00000110000100111100000000110000;
   assign mem[6084] = 32'b00000111111001000111110010100000;
   assign mem[6085] = 32'b11111100111001000001110110111000;
   assign mem[6086] = 32'b00000000000100100000001111101101;
   assign mem[6087] = 32'b00001111001110101000110000110000;
   assign mem[6088] = 32'b11111010100010101000110111001000;
   assign mem[6089] = 32'b11111001100100100010100111110000;
   assign mem[6090] = 32'b00000011110000011001000110010000;
   assign mem[6091] = 32'b00001001010110100010000100100000;
   assign mem[6092] = 32'b00000011101011010111001101110000;
   assign mem[6093] = 32'b11110001111100101011000100110000;
   assign mem[6094] = 32'b00000110011001111100011001110000;
   assign mem[6095] = 32'b11111000100001111000111010010000;
   assign mem[6096] = 32'b11111001011011010111101111010000;
   assign mem[6097] = 32'b11110111110111111000111001010000;
   assign mem[6098] = 32'b00000010101010100010111111011000;
   assign mem[6099] = 32'b11110110010100001111001000010000;
   assign mem[6100] = 32'b00000010111011000100110101100100;
   assign mem[6101] = 32'b11111111011111010101101010011101;
   assign mem[6102] = 32'b11111000001010110010110100011000;
   assign mem[6103] = 32'b11111101000111000001110100010000;
   assign mem[6104] = 32'b11111110001111000111011100110010;
   assign mem[6105] = 32'b00001000101101100111000010000000;
   assign mem[6106] = 32'b11111110010000111011001100011000;
   assign mem[6107] = 32'b11110111100011100000100000010000;
   assign mem[6108] = 32'b00000110001100010001001010011000;
   assign mem[6109] = 32'b00000000100001110010100100010010;
   assign mem[6110] = 32'b11110011110111011100100111000000;
   assign mem[6111] = 32'b00000001110110001110101110110000;
   assign mem[6112] = 32'b11111110010010011100010100010010;
   assign mem[6113] = 32'b00000001111110100111111110010110;
   assign mem[6114] = 32'b00000000100001001111000111011011;
   assign mem[6115] = 32'b11111110011011000110010101100010;
   assign mem[6116] = 32'b11111100010011111001010110110000;
   assign mem[6117] = 32'b00000101101100011000101101100000;
   assign mem[6118] = 32'b00000001100101100111111010011000;
   assign mem[6119] = 32'b11111110110011100101110101011010;
   assign mem[6120] = 32'b00000010010001010010010111111100;
   assign mem[6121] = 32'b11110000000100010001110010110000;
   assign mem[6122] = 32'b00000000100000101000110111001110;
   assign mem[6123] = 32'b11111011000110000100100101010000;
   assign mem[6124] = 32'b11111100101110100010011101111000;
   assign mem[6125] = 32'b00000010111000010110101001011100;
   assign mem[6126] = 32'b00001010000001101100000011100000;
   assign mem[6127] = 32'b11111111010000100101011011110011;
   assign mem[6128] = 32'b11111110001000111001000100011110;
   assign mem[6129] = 32'b00000010011100111010000000000000;
   assign mem[6130] = 32'b00000011000110101000000011100000;
   assign mem[6131] = 32'b11111001011011100100010011001000;
   assign mem[6132] = 32'b11111101101001001111100100110000;
   assign mem[6133] = 32'b11111100000101100010111011111000;
   assign mem[6134] = 32'b11111001111000111001001100101000;
   assign mem[6135] = 32'b00000000111001111110111001011001;
   assign mem[6136] = 32'b00000011110100001110000101000000;
   assign mem[6137] = 32'b11111111010000011000000101011010;
   assign mem[6138] = 32'b00000011111001101100010100000100;
   assign mem[6139] = 32'b00000000100101010010110100110110;
   assign mem[6140] = 32'b11111111001110101000001000010111;
   assign mem[6141] = 32'b11111000000111110001110111101000;
   assign mem[6142] = 32'b11111110110010000101100101010000;
   assign mem[6143] = 32'b11111101101101000100000000101000;
   assign mem[6144] = 32'b00000101010110101000010110001000;
   assign mem[6145] = 32'b00001001000110011001000111110000;
   assign mem[6146] = 32'b11111110101000000100010100100100;
   assign mem[6147] = 32'b11111000110010101010100000001000;
   assign mem[6148] = 32'b11111100100110111101101001010000;
   assign mem[6149] = 32'b00000011110110101110110110011000;
   assign mem[6150] = 32'b00000000100110011000000011001111;
   assign mem[6151] = 32'b11110100010111110010101110110000;
   assign mem[6152] = 32'b11111100010000001001110001011000;
   assign mem[6153] = 32'b11100111001101001101001000100000;
   assign mem[6154] = 32'b11110101011000101010111100100000;
   assign mem[6155] = 32'b00001100001101010110010101100000;
   assign mem[6156] = 32'b00001100101111001011101001100000;
   assign mem[6157] = 32'b11110110111110010000011001110000;
   assign mem[6158] = 32'b00000001101000001111001010010000;
   assign mem[6159] = 32'b11111000011111101100101100011000;
   assign mem[6160] = 32'b00001101110000010010000111010000;
   assign mem[6161] = 32'b11110101011000001110111101100000;
   assign mem[6162] = 32'b00000001111110011001001001000000;
   assign mem[6163] = 32'b11111100001110100010010101110100;
   assign mem[6164] = 32'b00000010010001010010001000001100;
   assign mem[6165] = 32'b11111010101010001111010011111000;
   assign mem[6166] = 32'b00000100001100100010000101111000;
   assign mem[6167] = 32'b00000001001110101000011010101100;
   assign mem[6168] = 32'b00000010001000101000100101000000;
   assign mem[6169] = 32'b11111111001110111110101101111100;
   assign mem[6170] = 32'b11110100010001110100011010100000;
   assign mem[6171] = 32'b11111110100111111110110110001110;
   assign mem[6172] = 32'b11101100100010110001011000100000;
   assign mem[6173] = 32'b11111100011011011000011111111000;
   assign mem[6174] = 32'b00000010001001100111111010111000;
   assign mem[6175] = 32'b00001001001001111000101110110000;
   assign mem[6176] = 32'b00000101000101111100101001010000;
   assign mem[6177] = 32'b00000001101110010100100101000010;
   assign mem[6178] = 32'b11111111101100000011000111111011;
   assign mem[6179] = 32'b11111111111110111101101010001010;
   assign mem[6180] = 32'b11111011100110110111100010110000;
   assign mem[6181] = 32'b11110111111011000011110010000000;
   assign mem[6182] = 32'b11110000001001100111100001100000;
   assign mem[6183] = 32'b11101000000001001000000001100000;
   assign mem[6184] = 32'b11110011100111100001100110100000;
   assign mem[6185] = 32'b00001010111101110101000111110000;
   assign mem[6186] = 32'b00010010111101110111111000000000;
   assign mem[6187] = 32'b11110110110111100101001101100000;
   assign mem[6188] = 32'b11110101000100011110001101000000;
   assign mem[6189] = 32'b11111001001000111010100001111000;
   assign mem[6190] = 32'b00000001110001000001000101101100;
   assign mem[6191] = 32'b11111101000000100001101001111100;
   assign mem[6192] = 32'b00000001001110101011011001111100;
   assign mem[6193] = 32'b00000011000011011110011111001000;
   assign mem[6194] = 32'b00000000101011000111001100101110;
   assign mem[6195] = 32'b11110000011011111000011001010000;
   assign mem[6196] = 32'b11111000111001000111001010100000;
   assign mem[6197] = 32'b00000001001010010111000001010110;
   assign mem[6198] = 32'b11111111100000100100100100110110;
   assign mem[6199] = 32'b00000001111011001111111010110100;
   assign mem[6200] = 32'b11111110101110000011101110010100;
   assign mem[6201] = 32'b00000011110111000101111100111100;
   assign mem[6202] = 32'b11110111101100110000100000010000;
   assign mem[6203] = 32'b00000011001100001010111101010000;
   assign mem[6204] = 32'b00000011010101000101111001000000;
   assign mem[6205] = 32'b11111111000110110000011101000101;
   assign mem[6206] = 32'b11111111000111000100011011001111;
   assign mem[6207] = 32'b11111110011000011111000010110100;
   assign mem[6208] = 32'b11111011110100111111111001000000;
   assign mem[6209] = 32'b11111111010010100011111100110101;
   assign mem[6210] = 32'b00000101100110001010010011111000;
   assign mem[6211] = 32'b11111100010011100010100000001000;
   assign mem[6212] = 32'b00000001000100101011110101010110;
   assign mem[6213] = 32'b11111111100101010010010101101111;
   assign mem[6214] = 32'b11110010101001101110110001110000;
   assign mem[6215] = 32'b11110101001110000011101001100000;
   assign mem[6216] = 32'b00000000100101100101011111100111;
   assign mem[6217] = 32'b00000000111101000101101011010001;
   assign mem[6218] = 32'b00000100011101000110001000011000;
   assign mem[6219] = 32'b00000101110001101110001100000000;
   assign mem[6220] = 32'b00001001101011010001000110110000;
   assign mem[6221] = 32'b11101111001011100110111100000000;
   assign mem[6222] = 32'b00000101001000111001101001000000;
   assign mem[6223] = 32'b11110001101101100100101111000000;
   assign mem[6224] = 32'b11110111111011101010100010010000;
   assign mem[6225] = 32'b00000111011111110110110000010000;
   assign mem[6226] = 32'b11111110100000100000101101000110;
   assign mem[6227] = 32'b11110010110000001111000011000000;
   assign mem[6228] = 32'b00000100101101001101110101011000;
   assign mem[6229] = 32'b11111101101001010101001001101000;
   assign mem[6230] = 32'b00000001110000001111011011111000;
   assign mem[6231] = 32'b11111100011110111101110000011000;
   assign mem[6232] = 32'b11111110100100100010011001111010;
   assign mem[6233] = 32'b11111101000010101101000000000000;
   assign mem[6234] = 32'b11111100100100011010011011001100;
   assign mem[6235] = 32'b11111101010001101010000000000000;
   assign mem[6236] = 32'b11111100110101101110010001001000;
   assign mem[6237] = 32'b11111111011001110111110111010010;
   assign mem[6238] = 32'b11111110100010100000111001010000;
   assign mem[6239] = 32'b00000001001100101000000110010100;
   assign mem[6240] = 32'b11111110010100000100111010010000;
   assign mem[6241] = 32'b00000110100111101010000100111000;
   assign mem[6242] = 32'b11110011111010000111001100110000;
   assign mem[6243] = 32'b11111110011000101111110001000100;
   assign mem[6244] = 32'b00000001000011011111010010001100;
   assign mem[6245] = 32'b00001000101010011000001110110000;
   assign mem[6246] = 32'b11111001110000110010010101100000;
   assign mem[6247] = 32'b00000011110111101100011010001000;
   assign mem[6248] = 32'b11111101000101110010000001001000;
   assign mem[6249] = 32'b11111111100111001110011110000111;
   assign mem[6250] = 32'b11111000111101110100000110010000;
   assign mem[6251] = 32'b00000111001110001001010110110000;
   assign mem[6252] = 32'b11111100001000010100000111110000;
   assign mem[6253] = 32'b11110111010000100010011000010000;
   assign mem[6254] = 32'b00001000001110001101001110110000;
   assign mem[6255] = 32'b11111111011011100110100011101101;
   assign mem[6256] = 32'b00000110100010001111100101100000;
   assign mem[6257] = 32'b00000111001111000010001110001000;
   assign mem[6258] = 32'b00000100010101000000001110100000;
   assign mem[6259] = 32'b11101000111110001011101110100000;
   assign mem[6260] = 32'b11111111000110110100110000110001;
   assign mem[6261] = 32'b11111011111101100000010111011000;
   assign mem[6262] = 32'b00000110000101000011100110101000;
   assign mem[6263] = 32'b00001000101101000101000110010000;
   assign mem[6264] = 32'b00000010000110111001100001010000;
   assign mem[6265] = 32'b11101100101101100010111000000000;
   assign mem[6266] = 32'b11111001010001101111110001100000;
   assign mem[6267] = 32'b00000010011010110111011010000000;
   assign mem[6268] = 32'b00000101001010010001100110111000;
   assign mem[6269] = 32'b11111100111100111110101111001000;
   assign mem[6270] = 32'b00000100010100101110101111010000;
   assign mem[6271] = 32'b00000111001001001111001111010000;
   assign mem[6272] = 32'b00000010010001101101100111001100;
   assign mem[6273] = 32'b11111001111110010101001101001000;
   assign mem[6274] = 32'b00000000110010101010001111011101;
   assign mem[6275] = 32'b11101111010100010001111000000000;
   assign mem[6276] = 32'b00000000101010100010100011010011;
   assign mem[6277] = 32'b11111101110001111111010011110100;
   assign mem[6278] = 32'b00000011111010100110100001111100;
   assign mem[6279] = 32'b11110110001011000010000010010000;
   assign mem[6280] = 32'b00000011100110101110110100010100;
   assign mem[6281] = 32'b11111101101110111111001000011000;
   assign mem[6282] = 32'b11110101011010100100011110010000;
   assign mem[6283] = 32'b11110100000100110100001011100000;
   assign mem[6284] = 32'b11111010000010111001111111011000;
   assign mem[6285] = 32'b00001101011111011110100000110000;
   assign mem[6286] = 32'b00000010101111101110110001101000;
   assign mem[6287] = 32'b00000000011000001100000101110000;
   assign mem[6288] = 32'b00000100010011100001101111011000;
   assign mem[6289] = 32'b00000000111111000100011110011100;
   assign mem[6290] = 32'b11111110010011011000000110101110;
   assign mem[6291] = 32'b11110011001111101100011001110000;
   assign mem[6292] = 32'b11110111001100000011110100010000;
   assign mem[6293] = 32'b11111001101010001011100111101000;
   assign mem[6294] = 32'b11110111011010011011110111000000;
   assign mem[6295] = 32'b00001011100111011100011110110000;
   assign mem[6296] = 32'b11111100110110111110000111100100;
   assign mem[6297] = 32'b11111101011101100111101011000000;
   assign mem[6298] = 32'b00000110110100100111010000010000;
   assign mem[6299] = 32'b11111011001000011000101111110000;
   assign mem[6300] = 32'b11110111111011010010001111010000;
   assign mem[6301] = 32'b00000011000111110111110111101000;
   assign mem[6302] = 32'b11101111011001011010001111000000;
   assign mem[6303] = 32'b00000100000000110110101101000000;
   assign mem[6304] = 32'b00000010001000000110010010100100;
   assign mem[6305] = 32'b00001001100010100100010001100000;
   assign mem[6306] = 32'b11111111111011011110010100010010;
   assign mem[6307] = 32'b00000101100111110110011110001000;
   assign mem[6308] = 32'b00000011101101010100000011101100;
   assign mem[6309] = 32'b11111001010010010010111000110000;
   assign mem[6310] = 32'b11111101000011101100001111110100;
   assign mem[6311] = 32'b00000001100000111101011000111000;
   assign mem[6312] = 32'b00000000101000100101010001001001;
   assign mem[6313] = 32'b00000110000010000010000100001000;
   assign mem[6314] = 32'b11111111011101001111101110100010;
   assign mem[6315] = 32'b11110000101001111011110011010000;
   assign mem[6316] = 32'b11111000101111010100110101100000;
   assign mem[6317] = 32'b00000011001010000011111001011100;
   assign mem[6318] = 32'b00000100101101100101000011000000;
   assign mem[6319] = 32'b11111011000000100101010000100000;
   assign mem[6320] = 32'b00000010011101111110110100101100;
   assign mem[6321] = 32'b00000000001100011101111100101111;
   assign mem[6322] = 32'b00000001011000001101111000110110;
   assign mem[6323] = 32'b00000101101111010001110001010000;
   assign mem[6324] = 32'b11111100111100000100110011001100;
   assign mem[6325] = 32'b11110000101010100100100100010000;
   assign mem[6326] = 32'b11110000110110011011010110110000;
   assign mem[6327] = 32'b00000011101000101010000100101000;
   assign mem[6328] = 32'b00000001001110010001111000111100;
   assign mem[6329] = 32'b00000010000101100101000110100100;
   assign mem[6330] = 32'b00001010100011110101001010100000;
   assign mem[6331] = 32'b11101101000010011100011001000000;
   assign mem[6332] = 32'b11111111111110000110100110110101;
   assign mem[6333] = 32'b11111010010111111101110110001000;
   assign mem[6334] = 32'b11100101101000010100011010100000;
   assign mem[6335] = 32'b00000000101110100100110000100000;
   assign mem[6336] = 32'b11111101111101001100110100010100;
   assign mem[6337] = 32'b11110111111000011000011011000000;
   assign mem[6338] = 32'b00000100110001001100001001011000;
   assign mem[6339] = 32'b00000101110100110001110100010000;
   assign mem[6340] = 32'b00000100011101001001100011111000;
   assign mem[6341] = 32'b11110001111011110000111011000000;
   assign mem[6342] = 32'b11111010001001000011110000110000;
   assign mem[6343] = 32'b11111110000100111111101001010110;
   assign mem[6344] = 32'b11111111111100100101010100111110;
   assign mem[6345] = 32'b11110100011010101101011011110000;
   assign mem[6346] = 32'b00000110100000011001101000011000;
   assign mem[6347] = 32'b00000010001110101000010101110000;
   assign mem[6348] = 32'b11111101101010100111000100111100;
   assign mem[6349] = 32'b11111110100110111110011011000100;
   assign mem[6350] = 32'b00000011000001011100100010101000;
   assign mem[6351] = 32'b11110111001110010111111110100000;
   assign mem[6352] = 32'b11111111110011000101010110110010;
   assign mem[6353] = 32'b00000001001001100010000010000110;
   assign mem[6354] = 32'b00000010000110110011010010101100;
   assign mem[6355] = 32'b11110010011101100101000011000000;
   assign mem[6356] = 32'b11111011010000001100011101110000;
   assign mem[6357] = 32'b00000011100010000101110011101100;
   assign mem[6358] = 32'b00000100100001101110110101101000;
   assign mem[6359] = 32'b00000100010111010001111011010000;
   assign mem[6360] = 32'b11110111101010011101010011100000;
   assign mem[6361] = 32'b11111110100111011011111001001000;
   assign mem[6362] = 32'b11111010010110011011111010111000;
   assign mem[6363] = 32'b11101110100011110101001101100000;
   assign mem[6364] = 32'b00000010111100100011011010111100;
   assign mem[6365] = 32'b00000001001110000111010011110110;
   assign mem[6366] = 32'b00000011110100101001000101010000;
   assign mem[6367] = 32'b00000100110010011011110011000000;
   assign mem[6368] = 32'b00000101101111101001010000101000;
   assign mem[6369] = 32'b11110011100010010111111100110000;
   assign mem[6370] = 32'b11110100010111110101110000010000;
   assign mem[6371] = 32'b00001001000111110011001011110000;
   assign mem[6372] = 32'b11111101011010100110000110111000;
   assign mem[6373] = 32'b11111000010111111001100000101000;
   assign mem[6374] = 32'b00001000010010001010000011110000;
   assign mem[6375] = 32'b00000000001101000001000110010001;
   assign mem[6376] = 32'b00000010110101111100011011111100;
   assign mem[6377] = 32'b00000101000101011111010011100000;
   assign mem[6378] = 32'b00000100011100010110110001110000;
   assign mem[6379] = 32'b11110001000001001111011011110000;
   assign mem[6380] = 32'b00000101001000101110010011100000;
   assign mem[6381] = 32'b00000110010110001000100011111000;
   assign mem[6382] = 32'b00000101010111100000001111001000;
   assign mem[6383] = 32'b11110100000110100111000000000000;
   assign mem[6384] = 32'b00001001110000010000000001100000;
   assign mem[6385] = 32'b11101111100110100000011111000000;
   assign mem[6386] = 32'b11110111101010100110011111000000;
   assign mem[6387] = 32'b11111000001001000001111100001000;
   assign mem[6388] = 32'b11111100001100110000100010100100;
   assign mem[6389] = 32'b11110100001111101101111100010000;
   assign mem[6390] = 32'b00000010010111001010100101001100;
   assign mem[6391] = 32'b00000001011111110100101100011110;
   assign mem[6392] = 32'b00001000001001001111000010000000;
   assign mem[6393] = 32'b11111100110101101101101100000100;
   assign mem[6394] = 32'b00000100101100110110100100100000;
   assign mem[6395] = 32'b11110110001000100110101101010000;
   assign mem[6396] = 32'b11110110001110010001001001000000;
   assign mem[6397] = 32'b11111111100100101110010111001000;
   assign mem[6398] = 32'b11111011111001111011000000011000;
   assign mem[6399] = 32'b11111011010101101011100010101000;
   assign mem[6400] = 32'b11110101001000000011100000100000;
   assign mem[6401] = 32'b00000100110110000001001110000000;
   assign mem[6402] = 32'b11111110100111111010000100001110;
   assign mem[6403] = 32'b00000000010011011000000100110000;
   assign mem[6404] = 32'b11111000010111010001111010101000;
   assign mem[6405] = 32'b00000010110010010101101000010000;
   assign mem[6406] = 32'b11111001010101100100011100101000;
   assign mem[6407] = 32'b11111100111100111101111001010000;
   assign mem[6408] = 32'b00000011111001001111011111010000;
   assign mem[6409] = 32'b00000001010110010011110001011000;
   assign mem[6410] = 32'b11110110000000010110010101010000;
   assign mem[6411] = 32'b11110110110110010101100111000000;
   assign mem[6412] = 32'b00000010011011001111110100101000;
   assign mem[6413] = 32'b00000110110000011011100101110000;
   assign mem[6414] = 32'b11111101110010111101010010111000;
   assign mem[6415] = 32'b00000101101101000100111011010000;
   assign mem[6416] = 32'b11111101110111101111011000100000;
   assign mem[6417] = 32'b00000011101110011010110110010000;
   assign mem[6418] = 32'b00000000010011101101000100011110;
   assign mem[6419] = 32'b11111111000011001000000011100011;
   assign mem[6420] = 32'b11111111101100010011011011010001;
   assign mem[6421] = 32'b11110101110010110110011010010000;
   assign mem[6422] = 32'b11110011100000010100101111110000;
   assign mem[6423] = 32'b11110010011110100010111001100000;
   assign mem[6424] = 32'b00000100100100101000011101001000;
   assign mem[6425] = 32'b11111000110010111011010001100000;
   assign mem[6426] = 32'b00000011001110001101010100011100;
   assign mem[6427] = 32'b11111000011010001001001011010000;
   assign mem[6428] = 32'b00001011110111001101110000100000;
   assign mem[6429] = 32'b00000011010111101111100000010100;
   assign mem[6430] = 32'b11110100101011110011010000110000;
   assign mem[6431] = 32'b11111110110001000100001101010100;
   assign mem[6432] = 32'b00000001111010101010001110111000;
   assign mem[6433] = 32'b00000000000011001001100000100100;
   assign mem[6434] = 32'b11111011001110111101101000111000;
   assign mem[6435] = 32'b11111101110110111100000000100000;
   assign mem[6436] = 32'b11101100110001000010100111000000;
   assign mem[6437] = 32'b00000110011101010011111001001000;
   assign mem[6438] = 32'b00000100111010000001110001001000;
   assign mem[6439] = 32'b11110010011001101001110010100000;
   assign mem[6440] = 32'b11111000111110000111011110111000;
   assign mem[6441] = 32'b00000101110000111100101011110000;
   assign mem[6442] = 32'b00001000010011010111111011100000;
   assign mem[6443] = 32'b00000101010110011100111111110000;
   assign mem[6444] = 32'b11110011000000000100110011100000;
   assign mem[6445] = 32'b00000010010100000110101000110000;
   assign mem[6446] = 32'b11110101110100111011100101100000;
   assign mem[6447] = 32'b00000100000001100001010001010000;
   assign mem[6448] = 32'b00000010000000101110110111101000;
   assign mem[6449] = 32'b11111100000001000111010111011000;
   assign mem[6450] = 32'b00000011111100100111011111110100;
   assign mem[6451] = 32'b00000101001011110110011000101000;
   assign mem[6452] = 32'b11110101101010011101001100010000;
   assign mem[6453] = 32'b11110110000111000101101000010000;
   assign mem[6454] = 32'b11111101101101000110011101000000;
   assign mem[6455] = 32'b11111010100110111111101100011000;
   assign mem[6456] = 32'b00001000011100011101011011000000;
   assign mem[6457] = 32'b11110111100100111111110100010000;
   assign mem[6458] = 32'b00000111000110110101110010111000;
   assign mem[6459] = 32'b00000100000101001111111010000000;
   assign mem[6460] = 32'b11111101011111110010000101010100;
   assign mem[6461] = 32'b00000011101111010011000000101000;
   assign mem[6462] = 32'b00000000111101101111011111101110;
   assign mem[6463] = 32'b00000010101011100011010110011000;
   assign mem[6464] = 32'b11111000100001100110000101101000;
   assign mem[6465] = 32'b11111111101111101111100010111001;
   assign mem[6466] = 32'b00000001101001101101110110011010;
   assign mem[6467] = 32'b11110111110010101010011000110000;
   assign mem[6468] = 32'b11111101110011100001010010001100;
   assign mem[6469] = 32'b00000011010011110010000010011000;
   assign mem[6470] = 32'b11111101111000010101110000111100;
   assign mem[6471] = 32'b00000100111110000110001100000000;
   assign mem[6472] = 32'b00000000111010111111011001111101;
   assign mem[6473] = 32'b00000111000100000011011111110000;
   assign mem[6474] = 32'b11110011010011111001010011110000;
   assign mem[6475] = 32'b11110110110101010110010001100000;
   assign mem[6476] = 32'b00000110011110110111010101001000;
   assign mem[6477] = 32'b00000001111000111100101011111100;
   assign mem[6478] = 32'b11110011111011110011010001110000;
   assign mem[6479] = 32'b00000001101011011101110111001100;
   assign mem[6480] = 32'b11111010110111110001110110110000;
   assign mem[6481] = 32'b11111001001011011110000011010000;
   assign mem[6482] = 32'b00001000101000001001111011000000;
   assign mem[6483] = 32'b00000111010010100010110101100000;
   assign mem[6484] = 32'b11111011001011011110001111101000;
   assign mem[6485] = 32'b00000001111100010011010010001010;
   assign mem[6486] = 32'b11110010000101111001010011010000;
   assign mem[6487] = 32'b00000111100110011010101001011000;
   assign mem[6488] = 32'b00000001110101110000110100100100;
   assign mem[6489] = 32'b11110011100110000010010100010000;
   assign mem[6490] = 32'b00000110001000010000000011111000;
   assign mem[6491] = 32'b11110110100110111011011001100000;
   assign mem[6492] = 32'b11111011110110101100100001000000;
   assign mem[6493] = 32'b11110110100101100111011010000000;
   assign mem[6494] = 32'b00000010110101001101101111000100;
   assign mem[6495] = 32'b11111111011111000011010011001100;
   assign mem[6496] = 32'b00001001101101110111000111100000;
   assign mem[6497] = 32'b00000011101011010101001011111100;
   assign mem[6498] = 32'b00000011010111110111110011001100;
   assign mem[6499] = 32'b00000010011000110001101111110000;
   assign mem[6500] = 32'b11111111110000011111000000111010;
   assign mem[6501] = 32'b00000010100111011001000101100000;
   assign mem[6502] = 32'b00000101001010111101101111110000;
   assign mem[6503] = 32'b11111110100010000001100100000010;
   assign mem[6504] = 32'b00000111011000011010111100001000;
   assign mem[6505] = 32'b11110010001100101001011101110000;
   assign mem[6506] = 32'b00000010000101111010111000000000;
   assign mem[6507] = 32'b00000101001111001100100101011000;
   assign mem[6508] = 32'b11111110000110100001100010110010;
   assign mem[6509] = 32'b11111011111110010010010110110000;
   assign mem[6510] = 32'b11111111011100111101010000101110;
   assign mem[6511] = 32'b11111001001101101100001110001000;
   assign mem[6512] = 32'b11111101110110101111100100001100;
   assign mem[6513] = 32'b11111001100111100100011100111000;
   assign mem[6514] = 32'b00000011100100001111110011000000;
   assign mem[6515] = 32'b11111111101111010110100010000111;
   assign mem[6516] = 32'b00000010100010010011001111010100;
   assign mem[6517] = 32'b11111001011101110100010001111000;
   assign mem[6518] = 32'b00000100010110001011101111011000;
   assign mem[6519] = 32'b00000110001001101101100001100000;
   assign mem[6520] = 32'b11111100010110011000101100001000;
   assign mem[6521] = 32'b11111101100010101000011000000100;
   assign mem[6522] = 32'b00001010001101010100010101100000;
   assign mem[6523] = 32'b11111001101111110111011111111000;
   assign mem[6524] = 32'b11110010010001001100011001010000;
   assign mem[6525] = 32'b00000010000111110110111001110100;
   assign mem[6526] = 32'b11111010010111111110010111100000;
   assign mem[6527] = 32'b11101111111000101011010000000000;
   assign mem[6528] = 32'b00001000011110110110010011010000;
   assign mem[6529] = 32'b11111110010101101011101000000100;
   assign mem[6530] = 32'b11110100111110100111010100100000;
   assign mem[6531] = 32'b11110100111110100000000000010000;
   assign mem[6532] = 32'b00000110010001001101110101010000;
   assign mem[6533] = 32'b00001001100010111011001000110000;
   assign mem[6534] = 32'b11111000011100011100000010011000;
   assign mem[6535] = 32'b00000100000101001110100110100000;
   assign mem[6536] = 32'b11110001100000100001011000000000;
   assign mem[6537] = 32'b00000001111000000001001100010100;
   assign mem[6538] = 32'b00000000010100111010010000010110;
   assign mem[6539] = 32'b11110111001101000010011111110000;
   assign mem[6540] = 32'b00000001011000010110101000111110;
   assign mem[6541] = 32'b11111001000111001101100101011000;
   assign mem[6542] = 32'b11111100011101111111110101010100;
   assign mem[6543] = 32'b11110011010011011011011110100000;
   assign mem[6544] = 32'b00000011001010100100010011001000;
   assign mem[6545] = 32'b00000001101101101110010001100100;
   assign mem[6546] = 32'b00000100101100100101101101101000;
   assign mem[6547] = 32'b11111000001010010001000110011000;
   assign mem[6548] = 32'b00000101101110001111000111000000;
   assign mem[6549] = 32'b00000110100101010000010011011000;
   assign mem[6550] = 32'b00000100101010000000000011011000;
   assign mem[6551] = 32'b11111101011000110100101001101100;
   assign mem[6552] = 32'b11111101111110100101111101001000;
   assign mem[6553] = 32'b11110011001110001100100010010000;
   assign mem[6554] = 32'b11111111000110111001011001100011;
   assign mem[6555] = 32'b11111111100111101011011110100000;
   assign mem[6556] = 32'b00000101010011010100011100111000;
   assign mem[6557] = 32'b11111111011011111001100111101111;
   assign mem[6558] = 32'b00000000000110101110010100011010;
   assign mem[6559] = 32'b00000011001110000101100011111100;
   assign mem[6560] = 32'b11111010110100101100010000100000;
   assign mem[6561] = 32'b11111010101110000110000100100000;
   assign mem[6562] = 32'b00000100101110000100011010111000;
   assign mem[6563] = 32'b00000101111010101110101000000000;
   assign mem[6564] = 32'b11111111010010110101011011000000;
   assign mem[6565] = 32'b00000010110110101111011010101100;
   assign mem[6566] = 32'b11101111010000111111100011100000;
   assign mem[6567] = 32'b00000101110010100011011101100000;
   assign mem[6568] = 32'b11111001001011001001000010111000;
   assign mem[6569] = 32'b11111001001000001100100110100000;
   assign mem[6570] = 32'b11111110110010101100001100111000;
   assign mem[6571] = 32'b11111110100011010101100001010010;
   assign mem[6572] = 32'b11110001101010010100010101000000;
   assign mem[6573] = 32'b11111010000100110010101100010000;
   assign mem[6574] = 32'b00000000100111100101001100001110;
   assign mem[6575] = 32'b11111010101100001111010110010000;
   assign mem[6576] = 32'b00000100110000101101001001110000;
   assign mem[6577] = 32'b00000000000100101111011000001110;
   assign mem[6578] = 32'b00000100010000001000001110001000;
   assign mem[6579] = 32'b00000010110101110111011000111100;
   assign mem[6580] = 32'b11111000110011001000010101011000;
   assign mem[6581] = 32'b11110111110000101001101100100000;
   assign mem[6582] = 32'b00000011010001011001010111001100;
   assign mem[6583] = 32'b00000110101000011111011011000000;
   assign mem[6584] = 32'b11111000011111100110001011100000;
   assign mem[6585] = 32'b11111001000100000100101000000000;
   assign mem[6586] = 32'b11110100010110101111101111010000;
   assign mem[6587] = 32'b00000010000000110011001011100000;
   assign mem[6588] = 32'b00000011100000000101100110100100;
   assign mem[6589] = 32'b11111000000100100001110011110000;
   assign mem[6590] = 32'b00000100111010110010001010001000;
   assign mem[6591] = 32'b11111000100110100000011101100000;
   assign mem[6592] = 32'b00001100010000111100101100010000;
   assign mem[6593] = 32'b00000011100001001010011001100000;
   assign mem[6594] = 32'b00000101101010100010001101110000;
   assign mem[6595] = 32'b11111000101111101010101000101000;
   assign mem[6596] = 32'b11111011000101101100101110011000;
   assign mem[6597] = 32'b11111011110001011011100000110000;
   assign mem[6598] = 32'b11111110111101000010100101010110;
   assign mem[6599] = 32'b11110100110001011011000100010000;
   assign mem[6600] = 32'b00000100111101000001100010101000;
   assign mem[6601] = 32'b00000001111110001001101111101110;
   assign mem[6602] = 32'b11110001100100000101100001100000;
   assign mem[6603] = 32'b11111001001010100001101001001000;
   assign mem[6604] = 32'b00000001100111010111111111101010;
   assign mem[6605] = 32'b11111111100100011110101100111001;
   assign mem[6606] = 32'b00000010100011000001011011101000;
   assign mem[6607] = 32'b00001000100111111111011001100000;
   assign mem[6608] = 32'b11111111111100001000110000011000;
   assign mem[6609] = 32'b00000100101001010000100001011000;
   assign mem[6610] = 32'b00000011010011110101010001010100;
   assign mem[6611] = 32'b11111101110111101011001100110100;
   assign mem[6612] = 32'b00001001001110010110000001000000;
   assign mem[6613] = 32'b00000001010000100110010011011110;
   assign mem[6614] = 32'b00000010011111110010101001111100;
   assign mem[6615] = 32'b11110010001100010000001110110000;
   assign mem[6616] = 32'b11110100000011011101011110110000;
   assign mem[6617] = 32'b00000111100010101110111011101000;
   assign mem[6618] = 32'b11111110110110010111001000010010;
   assign mem[6619] = 32'b11101110001111000111101001000000;
   assign mem[6620] = 32'b00000010011010010011100111111100;
   assign mem[6621] = 32'b00000010011101100011011010110100;
   assign mem[6622] = 32'b11111101000011000100010000000000;
   assign mem[6623] = 32'b11111000010100001101000110000000;
   assign mem[6624] = 32'b00000011010000100000010101000000;
   assign mem[6625] = 32'b11111100001000111111111111011100;
   assign mem[6626] = 32'b00000100001001010010000000001000;
   assign mem[6627] = 32'b11111111001101111011110001001111;
   assign mem[6628] = 32'b11110110100111011101100100000000;
   assign mem[6629] = 32'b00000100110101101101000100001000;
   assign mem[6630] = 32'b00000110011011111100111110001000;
   assign mem[6631] = 32'b11110111010011101111110101010000;
   assign mem[6632] = 32'b11101111110111111101100001000000;
   assign mem[6633] = 32'b11111001100011110110100110110000;
   assign mem[6634] = 32'b00000110110011011010010111111000;
   assign mem[6635] = 32'b11111111000100011110110010110000;
   assign mem[6636] = 32'b00000001111101100110100011000100;
   assign mem[6637] = 32'b11111101011101111100011001100100;
   assign mem[6638] = 32'b00000110010100001101101100011000;
   assign mem[6639] = 32'b00001001000100000111011110000000;
   assign mem[6640] = 32'b00000001011100011001101100100010;
   assign mem[6641] = 32'b11111001001111110011111100011000;
   assign mem[6642] = 32'b11111011101101011011111000100000;
   assign mem[6643] = 32'b11111001111100011100111010111000;
   assign mem[6644] = 32'b11111100011110100101100110101100;
   assign mem[6645] = 32'b00000000001100101011110100010111;
   assign mem[6646] = 32'b00000100011101110111010100101000;
   assign mem[6647] = 32'b11111011101010001011110001100000;
   assign mem[6648] = 32'b00000110001000000100010111101000;
   assign mem[6649] = 32'b00000111010101000101011101000000;
   assign mem[6650] = 32'b00000000000001110001101110011000;
   assign mem[6651] = 32'b00000100110100110001000010000000;
   assign mem[6652] = 32'b11111101011001111000101001010000;
   assign mem[6653] = 32'b00000010001100010000001000011000;
   assign mem[6654] = 32'b11111001110000101000010101111000;
   assign mem[6655] = 32'b11110101101000100000000001100000;
   assign mem[6656] = 32'b00001101010100000010000001010000;
   assign mem[6657] = 32'b11111011101011011010100110000000;
   assign mem[6658] = 32'b11110101010001110001001100010000;
   assign mem[6659] = 32'b00000100001001001011000011000000;
   assign mem[6660] = 32'b11111010000110010011111111001000;
   assign mem[6661] = 32'b00000100000110010111001101111000;
   assign mem[6662] = 32'b11101111101111110000010001000000;
   assign mem[6663] = 32'b00000101001010000111100011100000;
   assign mem[6664] = 32'b11110011101001101000110100110000;
   assign mem[6665] = 32'b11111110101001001000110111110010;
   assign mem[6666] = 32'b00000110001000100010000000000000;
   assign mem[6667] = 32'b11110110100011110001000111010000;
   assign mem[6668] = 32'b11111110101001001001110011101000;
   assign mem[6669] = 32'b00000100001100100111110010001000;
   assign mem[6670] = 32'b00000100001111101000100110110000;
   assign mem[6671] = 32'b11111011011000001100010001000000;
   assign mem[6672] = 32'b00000010110110101110011001100100;
   assign mem[6673] = 32'b11111001100100111111100011111000;
   assign mem[6674] = 32'b00000000011100100010101110011010;
   assign mem[6675] = 32'b00000001000011011001000111111010;
   assign mem[6676] = 32'b11111110101101111100101110000110;
   assign mem[6677] = 32'b11111010010110110011001010111000;
   assign mem[6678] = 32'b11111110100110100001100101111100;
   assign mem[6679] = 32'b11111010110001000100100111100000;
   assign mem[6680] = 32'b11111100111111001111001011100000;
   assign mem[6681] = 32'b00000001111101001101100000010100;
   assign mem[6682] = 32'b00000010000100010010101000001000;
   assign mem[6683] = 32'b11111010001101110001110110111000;
   assign mem[6684] = 32'b11111100101011010000010011100100;
   assign mem[6685] = 32'b11111100101100010011011100011000;
   assign mem[6686] = 32'b00000000011011111010001011111001;
   assign mem[6687] = 32'b00000010100111100111000111100100;
   assign mem[6688] = 32'b00000000111101011100100011110110;
   assign mem[6689] = 32'b00000100100111101100000100010000;
   assign mem[6690] = 32'b11111000100001110110101010001000;
   assign mem[6691] = 32'b11111001101100001111100001000000;
   assign mem[6692] = 32'b00001001100100010001111011000000;
   assign mem[6693] = 32'b00000011100111100110110110110100;
   assign mem[6694] = 32'b11111011110000010010010101101000;
   assign mem[6695] = 32'b11111111101111001111010001010101;
   assign mem[6696] = 32'b11110010001110100101011111110000;
   assign mem[6697] = 32'b00001001111111110100000100000000;
   assign mem[6698] = 32'b00000101101111001010011000100000;
   assign mem[6699] = 32'b11101110010110001111101001000000;
   assign mem[6700] = 32'b00000100111010000110000101011000;
   assign mem[6701] = 32'b00000001000100000101100110011010;
   assign mem[6702] = 32'b11101110000101111011010001100000;
   assign mem[6703] = 32'b00000110101100000010111010010000;
   assign mem[6704] = 32'b00001010001010000000010110000000;
   assign mem[6705] = 32'b11110000010100101001000110010000;
   assign mem[6706] = 32'b00000000011001111100000000011000;
   assign mem[6707] = 32'b00000100011101000110000100100000;
   assign mem[6708] = 32'b11111000101100111111111100101000;
   assign mem[6709] = 32'b11111110100111011111000011000000;
   assign mem[6710] = 32'b11110101101111111001101111100000;
   assign mem[6711] = 32'b11110101000000010001110011100000;
   assign mem[6712] = 32'b00000100111101010100111000011000;
   assign mem[6713] = 32'b00000100000100001101101010001000;
   assign mem[6714] = 32'b00000100110011011110101100110000;
   assign mem[6715] = 32'b00000001111010101010000010110010;
   assign mem[6716] = 32'b11110001100111111000111001010000;
   assign mem[6717] = 32'b00000011000111010010110111010000;
   assign mem[6718] = 32'b00000001001001011010110001101010;
   assign mem[6719] = 32'b11111111110010000000110010001001;
   assign mem[6720] = 32'b00000101000010010100110000000000;
   assign mem[6721] = 32'b11111100010001101101010111010100;
   assign mem[6722] = 32'b11111111100011011101000110100001;
   assign mem[6723] = 32'b11111011010101110000110011000000;
   assign mem[6724] = 32'b00000001000001100001100101000000;
   assign mem[6725] = 32'b11110001000001110011101000110000;
   assign mem[6726] = 32'b00001001110010111101101001110000;
   assign mem[6727] = 32'b00000001011010100011101110000100;
   assign mem[6728] = 32'b00000011001010110001010110101100;
   assign mem[6729] = 32'b00000011000100111111001110101000;
   assign mem[6730] = 32'b00000101101111100101001000001000;
   assign mem[6731] = 32'b00000011101100110111110100001100;
   assign mem[6732] = 32'b11110101000110011001011001010000;
   assign mem[6733] = 32'b11111011011111100101111111010000;
   assign mem[6734] = 32'b11111101101010100000001100000000;
   assign mem[6735] = 32'b11111000001001100001010111110000;
   assign mem[6736] = 32'b00000011110001110111101011011000;
   assign mem[6737] = 32'b11111111011111011101001110100010;
   assign mem[6738] = 32'b00000011000001110110110000000000;
   assign mem[6739] = 32'b00000100111001100011110110111000;
   assign mem[6740] = 32'b11110010110001101110010001100000;
   assign mem[6741] = 32'b11110111001010011101110000100000;
   assign mem[6742] = 32'b00000011011010010001001011000000;
   assign mem[6743] = 32'b11110100000001001101110011110000;
   assign mem[6744] = 32'b00000101011110000101011010000000;
   assign mem[6745] = 32'b00000000100000100000010001001000;
   assign mem[6746] = 32'b11111100100000001000000111110100;
   assign mem[6747] = 32'b11111011111001111001010111110000;
   assign mem[6748] = 32'b11111110110010101100101011010010;
   assign mem[6749] = 32'b00001000011001111000100100000000;
   assign mem[6750] = 32'b00000100000111000011111001010000;
   assign mem[6751] = 32'b11111010010111011010001110101000;
   assign mem[6752] = 32'b00000111001001000111011110001000;
   assign mem[6753] = 32'b11111000110100010011001000000000;
   assign mem[6754] = 32'b00000000111100100001101110010110;
   assign mem[6755] = 32'b00000010010110110100010001110000;
   assign mem[6756] = 32'b11111100100111110011111100000100;
   assign mem[6757] = 32'b11111000110000101101110100111000;
   assign mem[6758] = 32'b11111101110111110111011010110100;
   assign mem[6759] = 32'b11111110100111001000001001011100;
   assign mem[6760] = 32'b11101001011010000001010001100000;
   assign mem[6761] = 32'b11111110111000110111101000000100;
   assign mem[6762] = 32'b00000011110011011010110110011100;
   assign mem[6763] = 32'b00000111100101011001001110111000;
   assign mem[6764] = 32'b11110100100000110110100011000000;
   assign mem[6765] = 32'b00000011111011100100111001000100;
   assign mem[6766] = 32'b11101101111100010011111100000000;
   assign mem[6767] = 32'b00000010100110110000100010100100;
   assign mem[6768] = 32'b00000010111101110011110101101000;
   assign mem[6769] = 32'b11111110011000000100110100111100;
   assign mem[6770] = 32'b11111000001010010011011001111000;
   assign mem[6771] = 32'b11111101011111101011010110100100;
   assign mem[6772] = 32'b00000111000001111011111011110000;
   assign mem[6773] = 32'b00000111100110111000101010010000;
   assign mem[6774] = 32'b11111010000100000110110011110000;
   assign mem[6775] = 32'b11111011011111010111000001101000;
   assign mem[6776] = 32'b00000110011110000010100100101000;
   assign mem[6777] = 32'b00001000100010001100101000100000;
   assign mem[6778] = 32'b00000001111110100100001001111000;
   assign mem[6779] = 32'b11111110010001010110100100101110;
   assign mem[6780] = 32'b11111000001000001101110100100000;
   assign mem[6781] = 32'b00000000100011110111111110100110;
   assign mem[6782] = 32'b11111001000000001110001100111000;
   assign mem[6783] = 32'b11101111100010111100001110000000;
   assign mem[6784] = 32'b00001001001001101001001110110000;
   assign mem[6785] = 32'b00000001101001101011001101101000;
   assign mem[6786] = 32'b00000100010010001111101110010000;
   assign mem[6787] = 32'b11111100001101010111110100010100;
   assign mem[6788] = 32'b00000100000011000010101101110000;
   assign mem[6789] = 32'b00000010010111101001101101011000;
   assign mem[6790] = 32'b00000010011000101100001000000100;
   assign mem[6791] = 32'b11111010011101101111110110000000;
   assign mem[6792] = 32'b00001000110101110001111111010000;
   assign mem[6793] = 32'b00000100010101011010101000001000;
   assign mem[6794] = 32'b11111001010101100111111110100000;
   assign mem[6795] = 32'b11111011011011010001110001110000;
   assign mem[6796] = 32'b11111100011011111010110000010000;
   assign mem[6797] = 32'b11111101001011100010010100000100;
   assign mem[6798] = 32'b00000100001100110001110011100000;
   assign mem[6799] = 32'b11101110000100100001110011000000;
   assign mem[6800] = 32'b11111101110010110000001001111000;
   assign mem[6801] = 32'b11110111111100110101100001100000;
   assign mem[6802] = 32'b11111100101000100011110101100100;
   assign mem[6803] = 32'b11101101001100010011111111000000;
   assign mem[6804] = 32'b00000110001100111100110011111000;
   assign mem[6805] = 32'b00000001011010000100000111100100;
   assign mem[6806] = 32'b00000000011101011111011000111100;
   assign mem[6807] = 32'b11111001011101100011001101000000;
   assign mem[6808] = 32'b00000011100010000111001010001000;
   assign mem[6809] = 32'b00001001000010111101101010010000;
   assign mem[6810] = 32'b11111101001101001100000111001100;
   assign mem[6811] = 32'b00001000101111110000110111000000;
   assign mem[6812] = 32'b00000101001010101100110010001000;
   assign mem[6813] = 32'b00000011001101011000100101000100;
   assign mem[6814] = 32'b11110000100111100011001000110000;
   assign mem[6815] = 32'b11111110000100101000110010101110;
   assign mem[6816] = 32'b11111001001111001010101101001000;
   assign mem[6817] = 32'b00001001001101000100001101110000;
   assign mem[6818] = 32'b11111101001111000000100000100000;
   assign mem[6819] = 32'b11111001000010101011101111010000;
   assign mem[6820] = 32'b11110111001100001011000111100000;
   assign mem[6821] = 32'b00000100001111111000111110001000;
   assign mem[6822] = 32'b00000000011101110011001111010011;
   assign mem[6823] = 32'b00000011100011111100010011111100;
   assign mem[6824] = 32'b11111100001101110110010011001100;
   assign mem[6825] = 32'b11111111010100010011000010101011;
   assign mem[6826] = 32'b11101001011110110110100010100000;
   assign mem[6827] = 32'b00000001000110111100011110100010;
   assign mem[6828] = 32'b00000010011000001011011100001100;
   assign mem[6829] = 32'b11111101111010011101011101111000;
   assign mem[6830] = 32'b11111010010001001111001001110000;
   assign mem[6831] = 32'b00000010011000011110100000010100;
   assign mem[6832] = 32'b11111011000001010001110000000000;
   assign mem[6833] = 32'b00000001001100110100011000100100;
   assign mem[6834] = 32'b00000011111100001010010100110000;
   assign mem[6835] = 32'b11111110001100000010011010001100;
   assign mem[6836] = 32'b00000100001000110101110001111000;
   assign mem[6837] = 32'b00001000111001101110000000110000;
   assign mem[6838] = 32'b11111110111100011110001101101000;
   assign mem[6839] = 32'b00000010101101011110101001101100;
   assign mem[6840] = 32'b00000000010100001011111010100010;
   assign mem[6841] = 32'b11111000100100101100001001111000;
   assign mem[6842] = 32'b11110111111101100101110010100000;
   assign mem[6843] = 32'b11101111101101010101111111100000;
   assign mem[6844] = 32'b00001001111100011001010011000000;
   assign mem[6845] = 32'b00000010000010111110111001110100;
   assign mem[6846] = 32'b11111001010111010001100100111000;
   assign mem[6847] = 32'b11110011110010010001010100010000;
   assign mem[6848] = 32'b00000011011111000101110010111000;
   assign mem[6849] = 32'b00001001101011011101110000110000;
   assign mem[6850] = 32'b00000010100110111100001010111100;
   assign mem[6851] = 32'b11111011101110000110110011000000;
   assign mem[6852] = 32'b00000101000001001001110011111000;
   assign mem[6853] = 32'b11111110110011111011000101011010;
   assign mem[6854] = 32'b00000011000011011100010101101000;
   assign mem[6855] = 32'b11111100111101110010110001101000;
   assign mem[6856] = 32'b00000000011000100010001100111001;
   assign mem[6857] = 32'b00000100010001010100101010001000;
   assign mem[6858] = 32'b11111100111111000011110110101000;
   assign mem[6859] = 32'b00000000010010010001011001110100;
   assign mem[6860] = 32'b00000000001101111100010111011111;
   assign mem[6861] = 32'b11111010100101011010000001110000;
   assign mem[6862] = 32'b11111010001010101000011101010000;
   assign mem[6863] = 32'b11111010001110100000011100101000;
   assign mem[6864] = 32'b11111100111100001101110111111000;
   assign mem[6865] = 32'b00000011000011101100101000101100;
   assign mem[6866] = 32'b00000001101100000110000110110000;
   assign mem[6867] = 32'b00000110011110110110010111100000;
   assign mem[6868] = 32'b00000011010111010111011101100000;
   assign mem[6869] = 32'b00000001010101111001001011101110;
   assign mem[6870] = 32'b11111101110001101010101100100100;
   assign mem[6871] = 32'b11111011111010100000010010000000;
   assign mem[6872] = 32'b11111111010101111110110110001101;
   assign mem[6873] = 32'b00000001001001111010011001000100;
   assign mem[6874] = 32'b00000010011001100011011000000100;
   assign mem[6875] = 32'b00000001011110111100001011101010;
   assign mem[6876] = 32'b11111110101011011001111101000000;
   assign mem[6877] = 32'b11111111101000001101110110010111;
   assign mem[6878] = 32'b00000010010101100011011110100000;
   assign mem[6879] = 32'b00000001010110111001000000111100;
   assign mem[6880] = 32'b11110011101101011010011100100000;
   assign mem[6881] = 32'b11111101111000110110101010101000;
   assign mem[6882] = 32'b11110011100100010010110010000000;
   assign mem[6883] = 32'b11110101011111000101011001010000;
   assign mem[6884] = 32'b11111100111000101001100010011000;
   assign mem[6885] = 32'b11111101001100110101101100010100;
   assign mem[6886] = 32'b11111001011001100001101010101000;
   assign mem[6887] = 32'b00010001000010011000000101000000;
   assign mem[6888] = 32'b00000100010111010101101110101000;
   assign mem[6889] = 32'b11111110011111011100011001000110;
   assign mem[6890] = 32'b00001000000011101111000110110000;
   assign mem[6891] = 32'b11110100111111101101000101000000;
   assign mem[6892] = 32'b00000001111100101110101111100100;
   assign mem[6893] = 32'b11101111101110000110000111000000;
   assign mem[6894] = 32'b00000101001111110011001011011000;
   assign mem[6895] = 32'b11111001111101100110100001100000;
   assign mem[6896] = 32'b00000101111100111110000011010000;
   assign mem[6897] = 32'b11111111011000010000010010010111;
   assign mem[6898] = 32'b11111110100111000100011100110110;
   assign mem[6899] = 32'b00000100110000011100000010000000;
   assign mem[6900] = 32'b00000011001000100110110010010000;
   assign mem[6901] = 32'b00000001010110101110101110110000;
   assign mem[6902] = 32'b00000000101101101100011111100000;
   assign mem[6903] = 32'b11110111011101000000000011010000;
   assign mem[6904] = 32'b00000000001111101011111011000110;
   assign mem[6905] = 32'b11111010101000100110011000000000;
   assign mem[6906] = 32'b00000111100100100010000011100000;
   assign mem[6907] = 32'b11111110000011000100101100011100;
   assign mem[6908] = 32'b00000111010111101111010001101000;
   assign mem[6909] = 32'b00000100111111001100010001001000;
   assign mem[6910] = 32'b11111111111110010110111010001011;
   assign mem[6911] = 32'b11111101000011100111110111000000;
   assign mem[6912] = 32'b00000001111010101001110111100010;
   assign mem[6913] = 32'b11111111100000101110001011000011;
   assign mem[6914] = 32'b00000000100001111101110101100111;
   assign mem[6915] = 32'b11111111100100011110110011111001;
   assign mem[6916] = 32'b00000010001101100101000100001100;
   assign mem[6917] = 32'b11111100001111011000010011000100;
   assign mem[6918] = 32'b11111110110000101000101110101010;
   assign mem[6919] = 32'b11111010111000000011110011111000;
   assign mem[6920] = 32'b11110111111011011100100010000000;
   assign mem[6921] = 32'b11110110111101010110010101000000;
   assign mem[6922] = 32'b11111111001011000110000111011101;
   assign mem[6923] = 32'b11111111010000101011110101110100;
   assign mem[6924] = 32'b00000100000001110110110111110000;
   assign mem[6925] = 32'b00000110101111011100000101000000;
   assign mem[6926] = 32'b11111010010011001111101101011000;
   assign mem[6927] = 32'b11111101100110010001010011011000;
   assign mem[6928] = 32'b00000101000000101001000000111000;
   assign mem[6929] = 32'b11111110001100100111111111001110;
   assign mem[6930] = 32'b11111001001101010110011110001000;
   assign mem[6931] = 32'b11111110000010011001101111011100;
   assign mem[6932] = 32'b00000000100111101111110100011010;
   assign mem[6933] = 32'b11111101010001001011001000110100;
   assign mem[6934] = 32'b00000111001001010011111010000000;
   assign mem[6935] = 32'b11111011100100100100100111001000;
   assign mem[6936] = 32'b11110100111011011000011110100000;
   assign mem[6937] = 32'b00000010001101010001101110010100;
   assign mem[6938] = 32'b00001001110010110110100110000000;
   assign mem[6939] = 32'b00000001011101100001101100001100;
   assign mem[6940] = 32'b11111001100011101110000010101000;
   assign mem[6941] = 32'b11110111001000101101101100010000;
   assign mem[6942] = 32'b11111110001100010000110111101100;
   assign mem[6943] = 32'b11111110111000111010100110010110;
   assign mem[6944] = 32'b00000100100011000001110110101000;
   assign mem[6945] = 32'b00000111110001011111000101011000;
   assign mem[6946] = 32'b11110001000001100101110000110000;
   assign mem[6947] = 32'b00000001110110100101010001011100;
   assign mem[6948] = 32'b11111111000011110010110010011101;
   assign mem[6949] = 32'b00000111001111010011101100000000;
   assign mem[6950] = 32'b11111111001001010000000100110011;
   assign mem[6951] = 32'b00000100101110010100100000010000;
   assign mem[6952] = 32'b00000000001001110010001000001010;
   assign mem[6953] = 32'b11111100110001110110000000110000;
   assign mem[6954] = 32'b00000010110010011011101011011000;
   assign mem[6955] = 32'b11111110000000100101010001001010;
   assign mem[6956] = 32'b00000101010011001100100101010000;
   assign mem[6957] = 32'b11111100101000100111001011000000;
   assign mem[6958] = 32'b00000010011000011001000000000100;
   assign mem[6959] = 32'b00000100111100111110110000001000;
   assign mem[6960] = 32'b00000000101001100001000110010111;
   assign mem[6961] = 32'b11111110111101111001001100000000;
   assign mem[6962] = 32'b11111101101010100010100100001000;
   assign mem[6963] = 32'b11111110011101110100011001100010;
   assign mem[6964] = 32'b00000001111001101000110010010010;
   assign mem[6965] = 32'b00000000110000110001001010000011;
   assign mem[6966] = 32'b11111101101001101011001000010100;
   assign mem[6967] = 32'b00000110010001001001100101010000;
   assign mem[6968] = 32'b00000000011100111101100101010001;
   assign mem[6969] = 32'b00000010100100010010001100101100;
   assign mem[6970] = 32'b11110011111001011011110001110000;
   assign mem[6971] = 32'b00000001011010101001110110110110;
   assign mem[6972] = 32'b11111100100011001011101011111100;
   assign mem[6973] = 32'b11111101001111001000000011100000;
   assign mem[6974] = 32'b00000100010010111100101011110000;
   assign mem[6975] = 32'b00000011001000001110011001101100;
   assign mem[6976] = 32'b11111111010110111001010100011010;
   assign mem[6977] = 32'b00000000000000111011001000001000;
   assign mem[6978] = 32'b00000011001011000110110110111100;
   assign mem[6979] = 32'b00000111110110100100001000011000;
   assign mem[6980] = 32'b00000011011010011100110000011000;
   assign mem[6981] = 32'b11111001001111001101010100111000;
   assign mem[6982] = 32'b00001000011001000011101000010000;
   assign mem[6983] = 32'b11111111010010111010110001110001;
   assign mem[6984] = 32'b11111100010110001000101000111100;
   assign mem[6985] = 32'b11111101010011110011101111000100;
   assign mem[6986] = 32'b11111110011110010100011101110010;
   assign mem[6987] = 32'b11111110010101100110000100111000;
   assign mem[6988] = 32'b11111101100101011100010011100000;
   assign mem[6989] = 32'b11110110111001111100001101110000;
   assign mem[6990] = 32'b00000101001110000101100110010000;
   assign mem[6991] = 32'b11111110011111100101010110000100;
   assign mem[6992] = 32'b00000111111010110010110100101000;
   assign mem[6993] = 32'b11111111000100000100101011001101;
   assign mem[6994] = 32'b00000111100101110101001011000000;
   assign mem[6995] = 32'b11111001111001111100110110011000;
   assign mem[6996] = 32'b00000000001110101101101011111100;
   assign mem[6997] = 32'b00000001000010001110101010110000;
   assign mem[6998] = 32'b11111100111000010111110010001000;
   assign mem[6999] = 32'b11110011010101100101001101100000;
   assign mem[7000] = 32'b00000011110000001001100011100000;
   assign mem[7001] = 32'b11111100101011101010000001101100;
   assign mem[7002] = 32'b00001010001000110100100100010000;
   assign mem[7003] = 32'b00000001010000001011001110111000;
   assign mem[7004] = 32'b00000000101011100111111100110100;
   assign mem[7005] = 32'b11111110110111000111111101100000;
   assign mem[7006] = 32'b11111100011100110100011100010000;
   assign mem[7007] = 32'b11111101000011111011111011011100;
   assign mem[7008] = 32'b00000001110011110011111010001100;
   assign mem[7009] = 32'b11110110001000010001011100010000;
   assign mem[7010] = 32'b00000010011001011011000100010100;
   assign mem[7011] = 32'b11110011101111011101010110100000;
   assign mem[7012] = 32'b11111111011111010000110001011001;
   assign mem[7013] = 32'b11110011000001101110100010010000;
   assign mem[7014] = 32'b00000100010010101111001001010000;
   assign mem[7015] = 32'b11111001001000010101010111101000;
   assign mem[7016] = 32'b00000100010010011100000111100000;
   assign mem[7017] = 32'b00000011011000111001001101111000;
   assign mem[7018] = 32'b11111110110011000011010000111010;
   assign mem[7019] = 32'b00000100000001010001100011010000;
   assign mem[7020] = 32'b00000100001111010110010001011000;
   assign mem[7021] = 32'b11111001110001001111101010000000;
   assign mem[7022] = 32'b11111100111011010001000101100100;
   assign mem[7023] = 32'b11110011100101000001101110000000;
   assign mem[7024] = 32'b00000000001001101000100000110011;
   assign mem[7025] = 32'b00000001001111110101010001010100;
   assign mem[7026] = 32'b00000100101110100010010001001000;
   assign mem[7027] = 32'b11111111001010110100110000001110;
   assign mem[7028] = 32'b11111111000110000101011100010011;
   assign mem[7029] = 32'b11111111100000111100110101110111;
   assign mem[7030] = 32'b00000010101010110100110000111100;
   assign mem[7031] = 32'b11101111010101000111100011000000;
   assign mem[7032] = 32'b11110110010010001001000111100000;
   assign mem[7033] = 32'b11110110010110001011110111000000;
   assign mem[7034] = 32'b00000001011100010011101010010000;
   assign mem[7035] = 32'b11111100010111111001010101110100;
   assign mem[7036] = 32'b00000100100100100111111101000000;
   assign mem[7037] = 32'b11111110110011110001001100001110;
   assign mem[7038] = 32'b00000011001100101011010111001100;
   assign mem[7039] = 32'b00000010000110000000110111001000;
   assign mem[7040] = 32'b11111111101010110101110101100100;
   assign mem[7041] = 32'b11111010010111000000000101000000;
   assign mem[7042] = 32'b11111011100110001110001001111000;
   assign mem[7043] = 32'b00000000000100110001001000011001;
   assign mem[7044] = 32'b00000101010110101001010011100000;
   assign mem[7045] = 32'b00000011110000111000100101110100;
   assign mem[7046] = 32'b11101101010100001011110110100000;
   assign mem[7047] = 32'b11111011001011100001101110101000;
   assign mem[7048] = 32'b00000100110110011111111100000000;
   assign mem[7049] = 32'b00000101001111001000110110011000;
   assign mem[7050] = 32'b11111001110111010111001111011000;
   assign mem[7051] = 32'b11111001110001111011100001110000;
   assign mem[7052] = 32'b11111100111111000000001100011000;
   assign mem[7053] = 32'b00001110111100110000001011010000;
   assign mem[7054] = 32'b11110000111100010100011001100000;
   assign mem[7055] = 32'b00000111101111101110001111011000;
   assign mem[7056] = 32'b11111011100100110000100010010000;
   assign mem[7057] = 32'b11111000010111111010001000101000;
   assign mem[7058] = 32'b11111001000100001101000110110000;
   assign mem[7059] = 32'b00000101000010101101111110111000;
   assign mem[7060] = 32'b00000000011111000110011001111011;
   assign mem[7061] = 32'b11101000001010110100111100100000;
   assign mem[7062] = 32'b11110101000101011100010000000000;
   assign mem[7063] = 32'b11101110010100111110101000000000;
   assign mem[7064] = 32'b00000110000011101011101111110000;
   assign mem[7065] = 32'b11111111110001001001000110110011;
   assign mem[7066] = 32'b11111100000011100010110000101100;
   assign mem[7067] = 32'b11110110100100010010011010110000;
   assign mem[7068] = 32'b00001011100001100001100111000000;
   assign mem[7069] = 32'b00001000011111011001100011100000;
   assign mem[7070] = 32'b11101000001111100110000110100000;
   assign mem[7071] = 32'b11111101010101100110000011100000;
   assign mem[7072] = 32'b11111111011011011100111101000101;
   assign mem[7073] = 32'b00000000110101000011100011100010;
   assign mem[7074] = 32'b11111111101000010111000110111001;
   assign mem[7075] = 32'b00000011001111000010100000010000;
   assign mem[7076] = 32'b11100010101001111110011100100000;
   assign mem[7077] = 32'b00000010100010100010001010100000;
   assign mem[7078] = 32'b11111100111100111011000011111000;
   assign mem[7079] = 32'b00000010111001000101100110100100;
   assign mem[7080] = 32'b11111000001110110111001010101000;
   assign mem[7081] = 32'b00001001011000111011011111010000;
   assign mem[7082] = 32'b00000100011100111100110110100000;
   assign mem[7083] = 32'b00000001101000001010111110100100;
   assign mem[7084] = 32'b11110111110110101010000000000000;
   assign mem[7085] = 32'b00000010000101100000001011011000;
   assign mem[7086] = 32'b11110111011010110111001010110000;
   assign mem[7087] = 32'b00000111001100000010010000100000;
   assign mem[7088] = 32'b11110010110111100001000101010000;
   assign mem[7089] = 32'b11111001011100010000100110011000;
   assign mem[7090] = 32'b00000000001010100011111110100011;
   assign mem[7091] = 32'b11110010000010111010010110110000;
   assign mem[7092] = 32'b11111010111100011001100010110000;
   assign mem[7093] = 32'b11111010111000010011110111100000;
   assign mem[7094] = 32'b00000100101010101101110101011000;
   assign mem[7095] = 32'b00000010100011010001111001110100;
   assign mem[7096] = 32'b11111110001011110111111011100010;
   assign mem[7097] = 32'b11111010100111000100110001011000;
   assign mem[7098] = 32'b00000010100100000000100101111100;
   assign mem[7099] = 32'b00000000101100001111101100011100;
   assign mem[7100] = 32'b11111110100001100011110111111000;
   assign mem[7101] = 32'b00001001111101011000000010010000;
   assign mem[7102] = 32'b00000011100010111100001011010000;
   assign mem[7103] = 32'b00000111101111001111001000100000;
   assign mem[7104] = 32'b11110111011011100111100110110000;
   assign mem[7105] = 32'b11110011001111010111011000010000;
   assign mem[7106] = 32'b00001011101101100011111011110000;
   assign mem[7107] = 32'b00000000000110011101110110010010;
   assign mem[7108] = 32'b11110101010110000001010100100000;
   assign mem[7109] = 32'b11111011111111000001100100111000;
   assign mem[7110] = 32'b00000000111000010100111010111010;
   assign mem[7111] = 32'b00000100110111001110111011001000;
   assign mem[7112] = 32'b11111000100111101101101101000000;
   assign mem[7113] = 32'b00000111100010101001100001100000;
   assign mem[7114] = 32'b11111100101100000001010111110000;
   assign mem[7115] = 32'b11111010100001110001001011101000;
   assign mem[7116] = 32'b00000010011010010101011100110100;
   assign mem[7117] = 32'b00000100101011010001100001110000;
   assign mem[7118] = 32'b11111001101001010001000000101000;
   assign mem[7119] = 32'b11111010101101001110111001010000;
   assign mem[7120] = 32'b11101001110101110101001000000000;
   assign mem[7121] = 32'b11110110000000100101010011100000;
   assign mem[7122] = 32'b00001000010010000100110001010000;
   assign mem[7123] = 32'b00000010000100101001000011111100;
   assign mem[7124] = 32'b11110001101111110100101010000000;
   assign mem[7125] = 32'b11111111000001001100110101110010;
   assign mem[7126] = 32'b11111001011011001101011011011000;
   assign mem[7127] = 32'b00001101000110101110100101100000;
   assign mem[7128] = 32'b11111100111111100101100010110000;
   assign mem[7129] = 32'b00000001010111100001011111001000;
   assign mem[7130] = 32'b00000011000110001010100001010100;
   assign mem[7131] = 32'b00000000011001011010110010010011;
   assign mem[7132] = 32'b11111011100000111110101110000000;
   assign mem[7133] = 32'b11111010000100101011110110110000;
   assign mem[7134] = 32'b11111101111011101110101110111000;
   assign mem[7135] = 32'b00000010001011100101110001100000;
   assign mem[7136] = 32'b00000011101000010100111011111000;
   assign mem[7137] = 32'b11111110110100101000001111111110;
   assign mem[7138] = 32'b11111001110101100110111101110000;
   assign mem[7139] = 32'b11111111100101011110011010011011;
   assign mem[7140] = 32'b00000000110111010010011010101111;
   assign mem[7141] = 32'b00000000101010011011001000010011;
   assign mem[7142] = 32'b00000111000000011111101101001000;
   assign mem[7143] = 32'b11111111011001101101111010010110;
   assign mem[7144] = 32'b11111101110110111100111010110000;
   assign mem[7145] = 32'b11111001101011011100110101010000;
   assign mem[7146] = 32'b11111000100101010000110110110000;
   assign mem[7147] = 32'b00001000110001101101011010110000;
   assign mem[7148] = 32'b11111101000100000110110110001000;
   assign mem[7149] = 32'b11110111010101000111011100000000;
   assign mem[7150] = 32'b11110101100011101000100001110000;
   assign mem[7151] = 32'b11110110000000010010010000000000;
   assign mem[7152] = 32'b11100101111110110110001011000000;
   assign mem[7153] = 32'b11111100101111100000100110110000;
   assign mem[7154] = 32'b00000110011110011111000100110000;
   assign mem[7155] = 32'b11111111111000010101111101000100;
   assign mem[7156] = 32'b11110111101101000000100001010000;
   assign mem[7157] = 32'b11111110100000011110111101101100;
   assign mem[7158] = 32'b00000101101110100001001100010000;
   assign mem[7159] = 32'b00001001011101010110000000010000;
   assign mem[7160] = 32'b11110110111111100111011001100000;
   assign mem[7161] = 32'b11110000100101011111111011010000;
   assign mem[7162] = 32'b00000100010011110110100100011000;
   assign mem[7163] = 32'b11111000011010011101011000001000;
   assign mem[7164] = 32'b00000100010110010110100001000000;
   assign mem[7165] = 32'b11111111111100111000001110000110;
   assign mem[7166] = 32'b11111000110111101101111111110000;
   assign mem[7167] = 32'b11111001101101000110010111111000;
   assign mem[7168] = 32'b00000100011010001101110110010000;
   assign mem[7169] = 32'b00000100110111101000110000111000;
   assign mem[7170] = 32'b11111001000000011011001111000000;
   assign mem[7171] = 32'b11111011010101000111010010101000;
   assign mem[7172] = 32'b00000000000111011100110001010011;
   assign mem[7173] = 32'b11111011100001001101000101110000;
   assign mem[7174] = 32'b00000000100111110010010010011011;
   assign mem[7175] = 32'b11111011001011111100010000100000;
   assign mem[7176] = 32'b00000010101000101111001001010100;
   assign mem[7177] = 32'b11111110111001101010101011000110;
   assign mem[7178] = 32'b00001010001011100100101011110000;
   assign mem[7179] = 32'b11111101101010100101101110111100;
   assign mem[7180] = 32'b00000010100100000101100000110000;
   assign mem[7181] = 32'b11111000101001111100100010100000;
   assign mem[7182] = 32'b11111100001110110101000101001000;
   assign mem[7183] = 32'b11101111101011001010000010100000;
   assign mem[7184] = 32'b00000100110001100101111000100000;
   assign mem[7185] = 32'b00000110110001001001110010101000;
   assign mem[7186] = 32'b00000000001001100010111100111011;
   assign mem[7187] = 32'b11101111111000101000011101100000;
   assign mem[7188] = 32'b00001000101001110111110000000000;
   assign mem[7189] = 32'b00000111000001011001010101110000;
   assign mem[7190] = 32'b00000101011001111010001110110000;
   assign mem[7191] = 32'b00000001100011111001000101101110;
   assign mem[7192] = 32'b11111110001111110111111101111100;
   assign mem[7193] = 32'b11111111001010000101010110111111;
   assign mem[7194] = 32'b00000010111011111000110000100100;
   assign mem[7195] = 32'b00000010001001011000010011101100;
   assign mem[7196] = 32'b11111110011011100100101011011010;
   assign mem[7197] = 32'b11111111001010011101000100000000;
   assign mem[7198] = 32'b00000011100000001011111101010000;
   assign mem[7199] = 32'b11111110010000001000111100010000;
   assign mem[7200] = 32'b11110110010001100101001000000000;
   assign mem[7201] = 32'b00000001001101001110011001001100;
   assign mem[7202] = 32'b00000000101110000111110101000010;
   assign mem[7203] = 32'b11111111101110001111010011010100;
   assign mem[7204] = 32'b11111111111100110100100100111001;
   assign mem[7205] = 32'b00000011010000000111101110000000;
   assign mem[7206] = 32'b11110101100100000001000111010000;
   assign mem[7207] = 32'b00000111111100000110110000011000;
   assign mem[7208] = 32'b11110111000001011100110001000000;
   assign mem[7209] = 32'b11111111001000011011111110001111;
   assign mem[7210] = 32'b11111100100111001111111101111000;
   assign mem[7211] = 32'b11111001111011001011100110100000;
   assign mem[7212] = 32'b11111000100100101100110101010000;
   assign mem[7213] = 32'b11111000000110011111100000010000;
   assign mem[7214] = 32'b00000100101100000011011001100000;
   assign mem[7215] = 32'b00000000110101000010010110100011;
   assign mem[7216] = 32'b00000101011000010011010010111000;
   assign mem[7217] = 32'b00000000111010001100010110110100;
   assign mem[7218] = 32'b00000011110111011011101000011100;
   assign mem[7219] = 32'b00000011101100101110111110111000;
   assign mem[7220] = 32'b00000000010011100010011111101101;
   assign mem[7221] = 32'b00000010111111101011110111101000;
   assign mem[7222] = 32'b11111101000010100110100011111100;
   assign mem[7223] = 32'b11111101100010010010111110010000;
   assign mem[7224] = 32'b00000101110101100111101010100000;
   assign mem[7225] = 32'b00000010110110111010011010000100;
   assign mem[7226] = 32'b00000000101010000100110101001101;
   assign mem[7227] = 32'b11111111001001001010010010111011;
   assign mem[7228] = 32'b11110100011001001000010100010000;
   assign mem[7229] = 32'b00000100110100101100001010100000;
   assign mem[7230] = 32'b00000001101001011011001111001000;
   assign mem[7231] = 32'b00000010001101111011010111010100;
   assign mem[7232] = 32'b00000111111101000000110000000000;
   assign mem[7233] = 32'b11111100010001000001111100011100;
   assign mem[7234] = 32'b11111010101010011001001011110000;
   assign mem[7235] = 32'b11111000011101000011001000111000;
   assign mem[7236] = 32'b11111011001111100011001001111000;
   assign mem[7237] = 32'b00000001000000101000111100010000;
   assign mem[7238] = 32'b00000101110011001111011000000000;
   assign mem[7239] = 32'b11111000111000010101110011101000;
   assign mem[7240] = 32'b00000010010010011000101001000100;
   assign mem[7241] = 32'b11111111011110101011011010101010;
   assign mem[7242] = 32'b11111010011110101010011110000000;
   assign mem[7243] = 32'b11110100011101110101111011110000;
   assign mem[7244] = 32'b00000011010010110001000101111000;
   assign mem[7245] = 32'b00000001111011101111001101000000;
   assign mem[7246] = 32'b00000010010000101001100101111100;
   assign mem[7247] = 32'b00000100001010000011111000110000;
   assign mem[7248] = 32'b00000010011010101010100100010000;
   assign mem[7249] = 32'b00000010100111000101100111101100;
   assign mem[7250] = 32'b11111011101010100010110100101000;
   assign mem[7251] = 32'b11111010001011110010000011011000;
   assign mem[7252] = 32'b00001001011011100000101000010000;
   assign mem[7253] = 32'b11111101000100001000101110111100;
   assign mem[7254] = 32'b11111001101000111111110111010000;
   assign mem[7255] = 32'b11111001010110010010100000011000;
   assign mem[7256] = 32'b11111011110110001111001101110000;
   assign mem[7257] = 32'b00000110001011111011111110010000;
   assign mem[7258] = 32'b00000010000100101010001010010000;
   assign mem[7259] = 32'b11111100111001101101001001100000;
   assign mem[7260] = 32'b11111110110000001101001011100110;
   assign mem[7261] = 32'b00000001101000011011010001110010;
   assign mem[7262] = 32'b11110111001011111001101111000000;
   assign mem[7263] = 32'b11111101010101111001001011010100;
   assign mem[7264] = 32'b00001010001010101100011100000000;
   assign mem[7265] = 32'b11110101010101011001000011010000;
   assign mem[7266] = 32'b11111101110011000110101100001100;
   assign mem[7267] = 32'b11111111000111111000111011110111;
   assign mem[7268] = 32'b00000011001100000100011101011000;
   assign mem[7269] = 32'b00000001000000111110010100001100;
   assign mem[7270] = 32'b00000001011001100111000110110100;
   assign mem[7271] = 32'b11101001000011110011110100100000;
   assign mem[7272] = 32'b11101000011001010110100011000000;
   assign mem[7273] = 32'b11111000011011000011001001100000;
   assign mem[7274] = 32'b00000011111111011100011100100000;
   assign mem[7275] = 32'b00000011100010101010000011110000;
   assign mem[7276] = 32'b00000001100110011110111111100110;
   assign mem[7277] = 32'b11111010100010001011001011010000;
   assign mem[7278] = 32'b00000101101000111110011111101000;
   assign mem[7279] = 32'b00001001000111111000101100100000;
   assign mem[7280] = 32'b00000010000111110010111100000100;
   assign mem[7281] = 32'b11100101010100000100010110100000;
   assign mem[7282] = 32'b11101111110101111101110001100000;
   assign mem[7283] = 32'b11111010100100111011010011110000;
   assign mem[7284] = 32'b00000110011001101111000101110000;
   assign mem[7285] = 32'b00000100001011111101001100000000;
   assign mem[7286] = 32'b00000001000101111011100011110100;
   assign mem[7287] = 32'b00000001100011110001101011110110;
   assign mem[7288] = 32'b00001000100111011110000111110000;
   assign mem[7289] = 32'b00000101000110111010001001000000;
   assign mem[7290] = 32'b11111111111011001000100101011100;
   assign mem[7291] = 32'b00000001101100101110001010110010;
   assign mem[7292] = 32'b11110110011101101011001110000000;
   assign mem[7293] = 32'b11111001100110101111001011000000;
   assign mem[7294] = 32'b00000101000010110000100001100000;
   assign mem[7295] = 32'b11110001000110000101011000010000;
   assign mem[7296] = 32'b00000110110001011000100110100000;
   assign mem[7297] = 32'b00001101111001010011101110000000;
   assign mem[7298] = 32'b11111011001100111100100110110000;
   assign mem[7299] = 32'b00000000110010000101111100011010;
   assign mem[7300] = 32'b00000011011111010110101101000000;
   assign mem[7301] = 32'b11111011000100111010100101100000;
   assign mem[7302] = 32'b11101010100001010100000110000000;
   assign mem[7303] = 32'b11111010001111101011000101010000;
   assign mem[7304] = 32'b00000001011111001110010011100110;
   assign mem[7305] = 32'b00000100001101000000101010100000;
   assign mem[7306] = 32'b00000000111010101101010100010111;
   assign mem[7307] = 32'b11111111011000010100001001101011;
   assign mem[7308] = 32'b00001001010101100000011101010000;
   assign mem[7309] = 32'b00000000111110011101010100000101;
   assign mem[7310] = 32'b00000011111100111000000001010000;
   assign mem[7311] = 32'b00000110100100100010011100110000;
   assign mem[7312] = 32'b00000100001011110010101000101000;
   assign mem[7313] = 32'b11111111000100111010111110001110;
   assign mem[7314] = 32'b00000011001011010111100111010000;
   assign mem[7315] = 32'b11111011110110000010000000000000;
   assign mem[7316] = 32'b00000111110000101001100000010000;
   assign mem[7317] = 32'b00000111000000101100011101110000;
   assign mem[7318] = 32'b11111101100000111101111100000000;
   assign mem[7319] = 32'b11111010100101010010000011010000;
   assign mem[7320] = 32'b11111100110111111100111011110000;
   assign mem[7321] = 32'b11111110111111101110111000100110;
   assign mem[7322] = 32'b00001001100110100000011010010000;
   assign mem[7323] = 32'b11110011001110000000010100110000;
   assign mem[7324] = 32'b00000000101110001111100000011101;
   assign mem[7325] = 32'b00000110000011100011100001001000;
   assign mem[7326] = 32'b11111110100110100001100000000000;
   assign mem[7327] = 32'b11110101001011101111101010000000;
   assign mem[7328] = 32'b00000101101110010101111001010000;
   assign mem[7329] = 32'b00000111000001001010100100011000;
   assign mem[7330] = 32'b11110001111111101111101000010000;
   assign mem[7331] = 32'b11110100010110010111011100110000;
   assign mem[7332] = 32'b00001001110000110101011000000000;
   assign mem[7333] = 32'b00000100010110100110100101001000;
   assign mem[7334] = 32'b11111001101101110010010110001000;
   assign mem[7335] = 32'b11110111100001011011011010100000;
   assign mem[7336] = 32'b11111111111011000001000110011111;
   assign mem[7337] = 32'b00001111101111110101001111100000;
   assign mem[7338] = 32'b11111011100100010110100101110000;
   assign mem[7339] = 32'b11110111000001101001101011010000;
   assign mem[7340] = 32'b00000011110010100010010000010100;
   assign mem[7341] = 32'b11101100101111111100011011100000;
   assign mem[7342] = 32'b11110011011111101100110011010000;
   assign mem[7343] = 32'b11111100101111011001011001111000;
   assign mem[7344] = 32'b11111111101101111001110110110100;
   assign mem[7345] = 32'b11111111100001000111110001000011;
   assign mem[7346] = 32'b00000100011101100110010001011000;
   assign mem[7347] = 32'b00001010101001001111101110010000;
   assign mem[7348] = 32'b00000000110001010110011000001010;
   assign mem[7349] = 32'b00000010010110000011101111011100;
   assign mem[7350] = 32'b11110010011010000001111000000000;
   assign mem[7351] = 32'b11111100110101000000010101001000;
   assign mem[7352] = 32'b11111101101111101101000001111100;
   assign mem[7353] = 32'b11111101101100111010100010010000;
   assign mem[7354] = 32'b00000110001011110010110001110000;
   assign mem[7355] = 32'b00000001111010111010101000110000;
   assign mem[7356] = 32'b11100100110110000110101001000000;
   assign mem[7357] = 32'b00000110101000001000110110011000;
   assign mem[7358] = 32'b11111100010011110010011000110100;
   assign mem[7359] = 32'b00000101010110100110001000100000;
   assign mem[7360] = 32'b00000000110010111100010101011100;
   assign mem[7361] = 32'b00000001101000111111100110101000;
   assign mem[7362] = 32'b11111010010111111100100011011000;
   assign mem[7363] = 32'b11111111000101101111100000010111;
   assign mem[7364] = 32'b00000010100111010001100000001000;
   assign mem[7365] = 32'b11111010111101101101111010101000;
   assign mem[7366] = 32'b00000000011010010111011101010111;
   assign mem[7367] = 32'b00000010111001011110101000101100;
   assign mem[7368] = 32'b11111100011010100011010111111100;
   assign mem[7369] = 32'b11111101011111100110010011000000;
   assign mem[7370] = 32'b00000100101111100100110010000000;
   assign mem[7371] = 32'b11111101110010011000001100110100;
   assign mem[7372] = 32'b11111100110101011101101100011000;
   assign mem[7373] = 32'b11111000010010010100100111110000;
   assign mem[7374] = 32'b00000011000110000101011001011000;
   assign mem[7375] = 32'b11111110100001100000000000111010;
   assign mem[7376] = 32'b00000010111000000000111000010100;
   assign mem[7377] = 32'b11111101101000010010001101001100;
   assign mem[7378] = 32'b11111101110111011011000101111000;
   assign mem[7379] = 32'b00000110111111000101000100000000;
   assign mem[7380] = 32'b11111010010111010101011111001000;
   assign mem[7381] = 32'b11110000100000101010111001000000;
   assign mem[7382] = 32'b00000001010011101000011011110100;
   assign mem[7383] = 32'b11110100111100011000010011000000;
   assign mem[7384] = 32'b00000111011010001111100001000000;
   assign mem[7385] = 32'b00000001101011101100101011011010;
   assign mem[7386] = 32'b11110111000111001000110001010000;
   assign mem[7387] = 32'b00000001100101000000110101111100;
   assign mem[7388] = 32'b00000101000010001011001000100000;
   assign mem[7389] = 32'b00001000011100101100010111110000;
   assign mem[7390] = 32'b11111001100001110011110110010000;
   assign mem[7391] = 32'b00000010000110011110011010101100;
   assign mem[7392] = 32'b00000100011101110111000111100000;
   assign mem[7393] = 32'b00001000011110110000000111000000;
   assign mem[7394] = 32'b11111100000011010011000111101000;
   assign mem[7395] = 32'b11101111010110000100111011100000;
   assign mem[7396] = 32'b00001011001000111011100111010000;
   assign mem[7397] = 32'b11111110111010010100011010111110;
   assign mem[7398] = 32'b11110010111001001111010100110000;
   assign mem[7399] = 32'b11111011110100000100100011001000;
   assign mem[7400] = 32'b11110110111000100000001110100000;
   assign mem[7401] = 32'b11111001001000001000000111011000;
   assign mem[7402] = 32'b00000010100101001010101111000000;
   assign mem[7403] = 32'b11111101101000011001101110101100;
   assign mem[7404] = 32'b00000011011110000101011001101100;
   assign mem[7405] = 32'b11111110011100111001001011000110;
   assign mem[7406] = 32'b11111011010010101111100000100000;
   assign mem[7407] = 32'b00000011100001110010100111011000;
   assign mem[7408] = 32'b11111100010010110001100000011000;
   assign mem[7409] = 32'b00000010100111100110111100001100;
   assign mem[7410] = 32'b00000011101010011100000111011100;
   assign mem[7411] = 32'b11111101010111010010101000010100;
   assign mem[7412] = 32'b00000001000001000011010100011010;
   assign mem[7413] = 32'b00000001010001111111010011101100;
   assign mem[7414] = 32'b11111101111010000101101011000000;
   assign mem[7415] = 32'b00000011100101111100110011010100;
   assign mem[7416] = 32'b11111110001001011011111111000110;
   assign mem[7417] = 32'b00000011000111101101110101000000;
   assign mem[7418] = 32'b11111100101011101110011101000000;
   assign mem[7419] = 32'b00000001110101111100010111011010;
   assign mem[7420] = 32'b00000011011111001000101000011100;
   assign mem[7421] = 32'b11101111111000111011110110100000;
   assign mem[7422] = 32'b11111001010001001011001110000000;
   assign mem[7423] = 32'b11110110111111101000000000000000;
   assign mem[7424] = 32'b00000110011011011011111001110000;
   assign mem[7425] = 32'b00001000101111101111110010000000;
   assign mem[7426] = 32'b00000110100110011011111001101000;
   assign mem[7427] = 32'b11111001000110001110101001011000;
   assign mem[7428] = 32'b00000011001010111110011111101100;
   assign mem[7429] = 32'b00001000010110010101111000110000;
   assign mem[7430] = 32'b11110101100010000000101100000000;
   assign mem[7431] = 32'b00000100010101011101110101010000;
   assign mem[7432] = 32'b00001001000000110001111100010000;
   assign mem[7433] = 32'b00000010001101100010000101100100;
   assign mem[7434] = 32'b11101111111001000110011101000000;
   assign mem[7435] = 32'b11111100100110101111110001010100;
   assign mem[7436] = 32'b11110010110100011100001010110000;
   assign mem[7437] = 32'b00001010011001010011101001000000;
   assign mem[7438] = 32'b11111010100101100101110100001000;
   assign mem[7439] = 32'b11110001101100000111001000010000;
   assign mem[7440] = 32'b00000000110111000110011001101110;
   assign mem[7441] = 32'b00000000100010110010100110101110;
   assign mem[7442] = 32'b11110011101100010000000011000000;
   assign mem[7443] = 32'b11110001100101110010010001000000;
   assign mem[7444] = 32'b00000100100100110001111110110000;
   assign mem[7445] = 32'b00000100110000010010100111000000;
   assign mem[7446] = 32'b11110110111110110000000010000000;
   assign mem[7447] = 32'b00000010011000111101000000110000;
   assign mem[7448] = 32'b00000111110010111101010001101000;
   assign mem[7449] = 32'b00001010000101011100011000110000;
   assign mem[7450] = 32'b11111010001000110101100100111000;
   assign mem[7451] = 32'b00000011011110000001101100001000;
   assign mem[7452] = 32'b00000101001111100101100000001000;
   assign mem[7453] = 32'b00000011101010011111001001010100;
   assign mem[7454] = 32'b11111001000111111111011110010000;
   assign mem[7455] = 32'b00000110101101101001100111111000;
   assign mem[7456] = 32'b11111000101111001100010111000000;
   assign mem[7457] = 32'b00001000000110111010010100000000;
   assign mem[7458] = 32'b11110001110011000111100011100000;
   assign mem[7459] = 32'b11110111011001001001000010110000;
   assign mem[7460] = 32'b11100101001110111101010001000000;
   assign mem[7461] = 32'b00000011000010010010000011000100;
   assign mem[7462] = 32'b00000011010001001011110001111100;
   assign mem[7463] = 32'b00000101110000110010101100001000;
   assign mem[7464] = 32'b00000101000011101010000100000000;
   assign mem[7465] = 32'b00000100110011001101000111001000;
   assign mem[7466] = 32'b11011011010101111100101111000000;
   assign mem[7467] = 32'b00000011100001110110010001100100;
   assign mem[7468] = 32'b11111010010000110101110000101000;
   assign mem[7469] = 32'b00000010001101101100101101101000;
   assign mem[7470] = 32'b00000010101011100101000111110000;
   assign mem[7471] = 32'b11111101101010001110101100001000;
   assign mem[7472] = 32'b11110001000000100100101010100000;
   assign mem[7473] = 32'b11111110100000010100010100011110;
   assign mem[7474] = 32'b00000101001000000111001101010000;
   assign mem[7475] = 32'b00000000110111011100111101001101;
   assign mem[7476] = 32'b00000110000011010101001100000000;
   assign mem[7477] = 32'b11111111001101101000001000100011;
   assign mem[7478] = 32'b11111101000011110101110111010100;
   assign mem[7479] = 32'b00000001101000011111111010111110;
   assign mem[7480] = 32'b00000010110100001010001001101100;
   assign mem[7481] = 32'b11101101111100010110001010000000;
   assign mem[7482] = 32'b11111101111000100101011011010100;
   assign mem[7483] = 32'b11110111010010000110100000110000;
   assign mem[7484] = 32'b00000101101101010011010100011000;
   assign mem[7485] = 32'b00000010110101100010100001101000;
   assign mem[7486] = 32'b00000100101001100000110011000000;
   assign mem[7487] = 32'b11110001001110101111001011010000;
   assign mem[7488] = 32'b00000111101011001110110011110000;
   assign mem[7489] = 32'b00000110110111010100111110010000;
   assign mem[7490] = 32'b00000011100011001100011101010000;
   assign mem[7491] = 32'b11111100000000000101001110011000;
   assign mem[7492] = 32'b11111010010100000110111010011000;
   assign mem[7493] = 32'b11111101100100001110100110011100;
   assign mem[7494] = 32'b11111111001000011100000111111110;
   assign mem[7495] = 32'b11111011010000010101100110010000;
   assign mem[7496] = 32'b00000011010010010110001011000000;
   assign mem[7497] = 32'b00000100011110111111111111111000;
   assign mem[7498] = 32'b00000011011101011100101101001100;
   assign mem[7499] = 32'b00000000011001111111110000010011;
   assign mem[7500] = 32'b00000011010101000110111000010100;
   assign mem[7501] = 32'b00000001000001011001101000011100;
   assign mem[7502] = 32'b11110111111100111101010110110000;
   assign mem[7503] = 32'b11110111010100011110100001010000;
   assign mem[7504] = 32'b11111110010011011001011111010100;
   assign mem[7505] = 32'b00000000100000111000101111000111;
   assign mem[7506] = 32'b00000000111111010100111111110000;
   assign mem[7507] = 32'b11111010110100101010010011100000;
   assign mem[7508] = 32'b00000100111011011001001011101000;
   assign mem[7509] = 32'b00000100110111101001010111010000;
   assign mem[7510] = 32'b00000001001110101110000111110110;
   assign mem[7511] = 32'b11111101110011001100101011010000;
   assign mem[7512] = 32'b11111111010110111001110010011100;
   assign mem[7513] = 32'b11111101011111111110010111111000;
   assign mem[7514] = 32'b11111100010001011001110111001000;
   assign mem[7515] = 32'b00000011101000011110001011101100;
   assign mem[7516] = 32'b11111100110010010000000010011000;
   assign mem[7517] = 32'b11111110100101110001100110101000;
   assign mem[7518] = 32'b11111101010101101110011101011100;
   assign mem[7519] = 32'b11111100010000000101111000110000;
   assign mem[7520] = 32'b00000011101110101010010110101000;
   assign mem[7521] = 32'b11111101001010100100100001000100;
   assign mem[7522] = 32'b00000110000100110010111000101000;
   assign mem[7523] = 32'b11101100011001101100110101000000;
   assign mem[7524] = 32'b00000100000000001011010000000000;
   assign mem[7525] = 32'b00000100101001011100111110110000;
   assign mem[7526] = 32'b00000000000010110001000110110010;
   assign mem[7527] = 32'b00000100000010100100010110100000;
   assign mem[7528] = 32'b11111100000111000101100001001000;
   assign mem[7529] = 32'b11111111110101101101001100110101;
   assign mem[7530] = 32'b00000100010010011001100101001000;
   assign mem[7531] = 32'b00000001101101101011101000100010;
   assign mem[7532] = 32'b00000011001001101101011101110000;
   assign mem[7533] = 32'b11111011001111010010110100100000;
   assign mem[7534] = 32'b00000101010010011111000001101000;
   assign mem[7535] = 32'b11111110011110101011111001111110;
   assign mem[7536] = 32'b00000100100101011010010000000000;
   assign mem[7537] = 32'b11111101101000001011011001110000;
   assign mem[7538] = 32'b00000000100111110101100000001110;
   assign mem[7539] = 32'b11111101001011010010101100101000;
   assign mem[7540] = 32'b00000101100110100001000001110000;
   assign mem[7541] = 32'b00000001000001101010100000110000;
   assign mem[7542] = 32'b00000010000101101011100011010000;
   assign mem[7543] = 32'b11110101011111001111111010100000;
   assign mem[7544] = 32'b00000001010110100110010010010100;
   assign mem[7545] = 32'b00000000111100010010011101011101;
   assign mem[7546] = 32'b11111010100010001110111000001000;
   assign mem[7547] = 32'b11111101110011000011000110001100;
   assign mem[7548] = 32'b00001000010111010001000110110000;
   assign mem[7549] = 32'b11111101000101010001001111001100;
   assign mem[7550] = 32'b11111011111000011000001010100000;
   assign mem[7551] = 32'b11111111011000101100100111001000;
   assign mem[7552] = 32'b00000000110011100010101100110111;
   assign mem[7553] = 32'b00000101000001000110110000010000;
   assign mem[7554] = 32'b11111110101101111011111010010000;
   assign mem[7555] = 32'b00000001110101100001010010100110;
   assign mem[7556] = 32'b11111100111001101110101011010100;
   assign mem[7557] = 32'b11111101101101001100010100000000;
   assign mem[7558] = 32'b00000001000000001111000000001000;
   assign mem[7559] = 32'b00000000111001111110000010001111;
   assign mem[7560] = 32'b11110110111101100011010110000000;
   assign mem[7561] = 32'b11110111000101001011000101010000;
   assign mem[7562] = 32'b00000010100111110000001010100100;
   assign mem[7563] = 32'b11111111110101100110100011110110;
   assign mem[7564] = 32'b00000100111010100101100111000000;
   assign mem[7565] = 32'b00000000101001110011010111111011;
   assign mem[7566] = 32'b11110110101000011001111000010000;
   assign mem[7567] = 32'b00000010110111000101101111101000;
   assign mem[7568] = 32'b11111011010001110010111011111000;
   assign mem[7569] = 32'b00000010100000110010101001101000;
   assign mem[7570] = 32'b11111010101100011100100101110000;
   assign mem[7571] = 32'b11110101000010101001101001010000;
   assign mem[7572] = 32'b00000011111001101001110001101100;
   assign mem[7573] = 32'b11110101101101001100010001000000;
   assign mem[7574] = 32'b00000100110110000011101010100000;
   assign mem[7575] = 32'b11111011101011001011011100111000;
   assign mem[7576] = 32'b11101100000011111000001111100000;
   assign mem[7577] = 32'b11111100000111010011001110000100;
   assign mem[7578] = 32'b00000010100001011101010011011100;
   assign mem[7579] = 32'b00000100011100001001101101010000;
   assign mem[7580] = 32'b11111010100111101011100011011000;
   assign mem[7581] = 32'b11111101000010001011100101011000;
   assign mem[7582] = 32'b11111010111110111101001110011000;
   assign mem[7583] = 32'b11111111001100001100100000010111;
   assign mem[7584] = 32'b00000110011011101011100000000000;
   assign mem[7585] = 32'b00000011100111111001001101100100;
   assign mem[7586] = 32'b11110101000001011011110101100000;
   assign mem[7587] = 32'b00000101110101110001100100000000;
   assign mem[7588] = 32'b11111000001011011000010011110000;
   assign mem[7589] = 32'b00000000100111000000000101000101;
   assign mem[7590] = 32'b11111100100101011000101010001100;
   assign mem[7591] = 32'b00000000010111000011000011110100;
   assign mem[7592] = 32'b11110010011111010010010010110000;
   assign mem[7593] = 32'b00010001000000010100000111100000;
   assign mem[7594] = 32'b11111100100110000000101001110100;
   assign mem[7595] = 32'b11111011011101010001111001000000;
   assign mem[7596] = 32'b00000011010001011001100010011100;
   assign mem[7597] = 32'b11111100111000011001101100111100;
   assign mem[7598] = 32'b11111011001101001000110010001000;
   assign mem[7599] = 32'b00000111010011110101111100101000;
   assign mem[7600] = 32'b00000100001101100000110000000000;
   assign mem[7601] = 32'b11111101110101011110100000011100;
   assign mem[7602] = 32'b11110101001101100111101111010000;
   assign mem[7603] = 32'b11111010111010100010010100101000;
   assign mem[7604] = 32'b00001000110111001111001111010000;
   assign mem[7605] = 32'b11111011110011100011110000000000;
   assign mem[7606] = 32'b00000001000010000110101100101010;
   assign mem[7607] = 32'b00001011000101011100100111000000;
   assign mem[7608] = 32'b11111011011000100100010010000000;
   assign mem[7609] = 32'b11111001100101100101111000001000;
   assign mem[7610] = 32'b11101010010110110011010010100000;
   assign mem[7611] = 32'b11111110111100011110111100101010;
   assign mem[7612] = 32'b11111000001101000101100000101000;
   assign mem[7613] = 32'b11111101011010010100010011110100;
   assign mem[7614] = 32'b00000101100100001001110110000000;
   assign mem[7615] = 32'b00000000011101000011001010100001;
   assign mem[7616] = 32'b11101000101110000010011010000000;
   assign mem[7617] = 32'b00000010010010001111111011001100;
   assign mem[7618] = 32'b00000101011100001101001011101000;
   assign mem[7619] = 32'b00000111110100000101100111100000;
   assign mem[7620] = 32'b11111000000010011101000010001000;
   assign mem[7621] = 32'b11110111001101100010011101100000;
   assign mem[7622] = 32'b00000100101101101001000001100000;
   assign mem[7623] = 32'b11111110010000000101001011011110;
   assign mem[7624] = 32'b11111101110011110010011011011000;
   assign mem[7625] = 32'b11111101011010011001011101110100;
   assign mem[7626] = 32'b11111110011110111101101101010110;
   assign mem[7627] = 32'b00000011010110000001111011100000;
   assign mem[7628] = 32'b00000000001111110000011000010111;
   assign mem[7629] = 32'b11111100001101101000000000000000;
   assign mem[7630] = 32'b00000000010111110000010011000101;
   assign mem[7631] = 32'b11111001000011110100000110100000;
   assign mem[7632] = 32'b00000001100011101001010101010010;
   assign mem[7633] = 32'b11110111100011110011000010000000;
   assign mem[7634] = 32'b00000011101101110111110110010000;
   assign mem[7635] = 32'b11111111011011011011100111000111;
   assign mem[7636] = 32'b00000110001111010000001010010000;
   assign mem[7637] = 32'b00000100001000100010000001110000;
   assign mem[7638] = 32'b11111111101101001101000110010010;
   assign mem[7639] = 32'b11111111101110000010011111101010;
   assign mem[7640] = 32'b00000001110100001010011100000010;
   assign mem[7641] = 32'b00000101111110011101101100001000;
   assign mem[7642] = 32'b00000101010001000011101000100000;
   assign mem[7643] = 32'b00000100001100111011010111101000;
   assign mem[7644] = 32'b11111110110110010111011010000000;
   assign mem[7645] = 32'b11111011111111011000010000001000;
   assign mem[7646] = 32'b11111101101110110000001000110000;
   assign mem[7647] = 32'b00001100000101010011111010000000;
   assign mem[7648] = 32'b11111110111110000101010101101110;
   assign mem[7649] = 32'b11101101001001010110111110000000;
   assign mem[7650] = 32'b00000100001011100000100111000000;
   assign mem[7651] = 32'b11111101111001000110001100110000;
   assign mem[7652] = 32'b00000000111111011010010110000010;
   assign mem[7653] = 32'b11110100000010000001001111110000;
   assign mem[7654] = 32'b00000100100011111001110101110000;
   assign mem[7655] = 32'b11111110011011000000010000000110;
   assign mem[7656] = 32'b00000001111000011010110111010110;
   assign mem[7657] = 32'b11111101011101100001011010101100;
   assign mem[7658] = 32'b11111011011010010100000100000000;
   assign mem[7659] = 32'b00000011001000100010111000001000;
   assign mem[7660] = 32'b00000000011100110110001110110100;
   assign mem[7661] = 32'b00000001000010101001100101000000;
   assign mem[7662] = 32'b11111100001000011100010110100000;
   assign mem[7663] = 32'b11111011000000110110100101111000;
   assign mem[7664] = 32'b11111110111000010111001001001000;
   assign mem[7665] = 32'b00000011011110011110101001101000;
   assign mem[7666] = 32'b00000110011000010011000011110000;
   assign mem[7667] = 32'b00000000101100101100001010001111;
   assign mem[7668] = 32'b11111110101011100001110100111110;
   assign mem[7669] = 32'b00000001110111001110001010111010;
   assign mem[7670] = 32'b00000001100111011100010011010000;
   assign mem[7671] = 32'b00000001111111010000011010010010;
   assign mem[7672] = 32'b11111100110110100001011001101000;
   assign mem[7673] = 32'b11110010010000000000111010100000;
   assign mem[7674] = 32'b00000001011101000011010000011000;
   assign mem[7675] = 32'b00000011100111010010101101011000;
   assign mem[7676] = 32'b00000001100111011101100111100100;
   assign mem[7677] = 32'b11111100010100010011011111000000;
   assign mem[7678] = 32'b11111100001101101101010100111100;
   assign mem[7679] = 32'b00000100100000001111111100100000;
   assign mem[7680] = 32'b00001010001001000101010000000000;
   assign mem[7681] = 32'b11110101100100011001010000010000;
   assign mem[7682] = 32'b11111100001000101101000010011100;
   assign mem[7683] = 32'b00000000010100111111010111100101;
   assign mem[7684] = 32'b00000101010011010111001101000000;
   assign mem[7685] = 32'b11111101101010110011100110000100;
   assign mem[7686] = 32'b00000001010011011110101011111000;
   assign mem[7687] = 32'b11111011011111110101011110111000;
   assign mem[7688] = 32'b00000011101100010010000101001000;
   assign mem[7689] = 32'b00000000000111100001011110111111;
   assign mem[7690] = 32'b00001001000100101101011010110000;
   assign mem[7691] = 32'b00000011101001111001100101010100;
   assign mem[7692] = 32'b00000100110011001011001100101000;
   assign mem[7693] = 32'b11110110000110000010010101000000;
   assign mem[7694] = 32'b11111010001011010100100100101000;
   assign mem[7695] = 32'b00000111000100010111100000010000;
   assign mem[7696] = 32'b11111101011000101011111110000000;
   assign mem[7697] = 32'b00001101000010011011111110010000;
   assign mem[7698] = 32'b11111001110101111010100111001000;
   assign mem[7699] = 32'b11101010110100011010111110100000;
   assign mem[7700] = 32'b00000001101100111101110010111000;
   assign mem[7701] = 32'b11111110101100100100110101101110;
   assign mem[7702] = 32'b11111110100100100001110110000110;
   assign mem[7703] = 32'b00000000010110010001010001100111;
   assign mem[7704] = 32'b00001001111001100010001000010000;
   assign mem[7705] = 32'b00000000010110010011011111101010;
   assign mem[7706] = 32'b11111101001011101001001010001000;
   assign mem[7707] = 32'b11110011110111110110101111100000;
   assign mem[7708] = 32'b00000010111110001000111111111000;
   assign mem[7709] = 32'b11111111000001111100110010100110;
   assign mem[7710] = 32'b11110100010100001111000000010000;
   assign mem[7711] = 32'b11110000000000110000101111100000;
   assign mem[7712] = 32'b11111111101100101000010000110100;
   assign mem[7713] = 32'b11111111111111000101001001001000;
   assign mem[7714] = 32'b11111110010001101110011110010010;
   assign mem[7715] = 32'b00000001111000100011100001110000;
   assign mem[7716] = 32'b11110101011100001111110000110000;
   assign mem[7717] = 32'b00000000000101110101001010000100;
   assign mem[7718] = 32'b11111001111011011101101110101000;
   assign mem[7719] = 32'b00000111011110001101111111001000;
   assign mem[7720] = 32'b11111101011110011111100000101100;
   assign mem[7721] = 32'b00000010000010100010100011001000;
   assign mem[7722] = 32'b00000100000001001111011111011000;
   assign mem[7723] = 32'b00000001101110101010001101110010;
   assign mem[7724] = 32'b11111101100001110101110001010000;
   assign mem[7725] = 32'b00000010010100010001101001001000;
   assign mem[7726] = 32'b11111101000100001110100111110100;
   assign mem[7727] = 32'b00000011001010001001011111011100;
   assign mem[7728] = 32'b11110001011111001100001101110000;
   assign mem[7729] = 32'b11111100100100110100010010010000;
   assign mem[7730] = 32'b11111110111010011100011001101010;
   assign mem[7731] = 32'b11111110100110101000000001010110;
   assign mem[7732] = 32'b11111010011000111101101001111000;
   assign mem[7733] = 32'b11111101011010111001110100011000;
   assign mem[7734] = 32'b00000011011001000111100110110100;
   assign mem[7735] = 32'b00000000010101000000111001010011;
   assign mem[7736] = 32'b00000100011100100101101101100000;
   assign mem[7737] = 32'b00000000101001010100110101011000;
   assign mem[7738] = 32'b00000001010001010001000000111100;
   assign mem[7739] = 32'b11111110010110101111000111010110;
   assign mem[7740] = 32'b00000011110001011110111100101000;
   assign mem[7741] = 32'b00000001011001110110110001001000;
   assign mem[7742] = 32'b11111011111101111111000011100000;
   assign mem[7743] = 32'b11110111010100110010110011010000;
   assign mem[7744] = 32'b00000000001000001011010000000101;
   assign mem[7745] = 32'b00000001101001000100110111000110;
   assign mem[7746] = 32'b11111101111000011111010111011100;
   assign mem[7747] = 32'b00001111000000000100111110000000;
   assign mem[7748] = 32'b11110011010010110100110110100000;
   assign mem[7749] = 32'b11111011110001110111001000101000;
   assign mem[7750] = 32'b00000100001000101110101000110000;
   assign mem[7751] = 32'b00000110100011100110001010000000;
   assign mem[7752] = 32'b11111101001001100111010100000000;
   assign mem[7753] = 32'b00000000110110010110010010010001;
   assign mem[7754] = 32'b11111101110101010000000011110000;
   assign mem[7755] = 32'b00000000100101111010000000001010;
   assign mem[7756] = 32'b00000101101100010100110010100000;
   assign mem[7757] = 32'b00000100110001010000101101001000;
   assign mem[7758] = 32'b00000000011001111011100010001100;
   assign mem[7759] = 32'b11111101100101111011100000100000;
   assign mem[7760] = 32'b11111111110101111011101010111011;
   assign mem[7761] = 32'b11110001010100110001111011100000;
   assign mem[7762] = 32'b00000111011100001011000101101000;
   assign mem[7763] = 32'b11111111110100010000100011010100;
   assign mem[7764] = 32'b11111100011001001100101000110100;
   assign mem[7765] = 32'b00000011110111100101001001100100;
   assign mem[7766] = 32'b11111001110111000001010011100000;
   assign mem[7767] = 32'b00001000010110010110101000110000;
   assign mem[7768] = 32'b11110110010101110001110110000000;
   assign mem[7769] = 32'b11110111101101111011011111100000;
   assign mem[7770] = 32'b11110010000101111111100000010000;
   assign mem[7771] = 32'b00000100111011100110001101010000;
   assign mem[7772] = 32'b00000100010100111001101100010000;
   assign mem[7773] = 32'b11111011011111010011011111000000;
   assign mem[7774] = 32'b11110001110001111011111100010000;
   assign mem[7775] = 32'b00000100100100101011110101000000;
   assign mem[7776] = 32'b11111111000011100100000001101101;
   assign mem[7777] = 32'b00001010000110110111001111100000;
   assign mem[7778] = 32'b11111101000100001110001011001100;
   assign mem[7779] = 32'b11111011101111110110100010101000;
   assign mem[7780] = 32'b11110010000101101111010011100000;
   assign mem[7781] = 32'b00000111010110010001001101101000;
   assign mem[7782] = 32'b00000101101001101101000010100000;
   assign mem[7783] = 32'b00000011001000010100111101110000;
   assign mem[7784] = 32'b00000001110010000101010100100110;
   assign mem[7785] = 32'b00000011111001111010100111000000;
   assign mem[7786] = 32'b00000010010010011101001101011000;
   assign mem[7787] = 32'b11111110001101011001111011111110;
   assign mem[7788] = 32'b11111101001001010101010010110000;
   assign mem[7789] = 32'b00000100010110000001100100010000;
   assign mem[7790] = 32'b11111100001001101101110100111000;
   assign mem[7791] = 32'b11111111100111111101100100001001;
   assign mem[7792] = 32'b11110101111111001100010110010000;
   assign mem[7793] = 32'b00000101000000000110101100111000;
   assign mem[7794] = 32'b00000100010011101111110100001000;
   assign mem[7795] = 32'b00000101000101001001100111000000;
   assign mem[7796] = 32'b11110100010110010111110000110000;
   assign mem[7797] = 32'b11111010011111110000110110101000;
   assign mem[7798] = 32'b00000011010100111001000000111100;
   assign mem[7799] = 32'b00000010011111001000101001111100;
   assign mem[7800] = 32'b11111010000111010111110010101000;
   assign mem[7801] = 32'b11100101001011011100100100100000;
   assign mem[7802] = 32'b00000101101000101100010000110000;
   assign mem[7803] = 32'b11111101001111000100100110001100;
   assign mem[7804] = 32'b00001001100110110110010100010000;
   assign mem[7805] = 32'b00000010010011001110110010111000;
   assign mem[7806] = 32'b00001000000101011000001101100000;
   assign mem[7807] = 32'b11101111110000100100110101000000;
   assign mem[7808] = 32'b00000001001000000011100010010100;
   assign mem[7809] = 32'b00000001010110011010010011111110;
   assign mem[7810] = 32'b11111101010010111011100101010100;
   assign mem[7811] = 32'b11110101100100101100111011100000;
   assign mem[7812] = 32'b00001011110010101101111110110000;
   assign mem[7813] = 32'b11111000010101110011110010001000;
   assign mem[7814] = 32'b00001000111001011001001001110000;
   assign mem[7815] = 32'b00001011010000001000110111010000;
   assign mem[7816] = 32'b00001010111010111111000100110000;
   assign mem[7817] = 32'b11110101101001110010010101000000;
   assign mem[7818] = 32'b11111010001010111101000110111000;
   assign mem[7819] = 32'b11110101101111000011001110010000;
   assign mem[7820] = 32'b11111000001100001011111011101000;
   assign mem[7821] = 32'b11110000001100001100111001000000;
   assign mem[7822] = 32'b11111011101100110110001000010000;
   assign mem[7823] = 32'b11111101010010011100000000110000;
   assign mem[7824] = 32'b00000101110001011011111100011000;
   assign mem[7825] = 32'b00000010010111000100101101101000;
   assign mem[7826] = 32'b00000000101100001111110110110110;
   assign mem[7827] = 32'b11101011000111110100101100000000;
   assign mem[7828] = 32'b00000101011101111101000011100000;
   assign mem[7829] = 32'b00000110110000111000011000111000;
   assign mem[7830] = 32'b11110011001010110011100111100000;
   assign mem[7831] = 32'b00000000100011000011010001100001;
   assign mem[7832] = 32'b00000000000001010110111001010101;
   assign mem[7833] = 32'b11111111110010011101111010010001;
   assign mem[7834] = 32'b11110101110000011101100111000000;
   assign mem[7835] = 32'b11111011001110000110111011010000;
   assign mem[7836] = 32'b11111111001110100110100001111010;
   assign mem[7837] = 32'b00000011001110101000100100000000;
   assign mem[7838] = 32'b00000100101011100010000010100000;
   assign mem[7839] = 32'b11111101100011010100110110100100;
   assign mem[7840] = 32'b11110111011010000001111010110000;
   assign mem[7841] = 32'b11101010100010111010000000100000;
   assign mem[7842] = 32'b11110100110011111101111000000000;
   assign mem[7843] = 32'b11111111011101111010110111100111;
   assign mem[7844] = 32'b00000000101100010000001111110101;
   assign mem[7845] = 32'b00000001100110111100101001111100;
   assign mem[7846] = 32'b00000000111000000100011010110001;
   assign mem[7847] = 32'b11111010111011011010111011001000;
   assign mem[7848] = 32'b11111111110010100000100011010010;
   assign mem[7849] = 32'b00001000001011010010001110010000;
   assign mem[7850] = 32'b11110100101111111001010011000000;
   assign mem[7851] = 32'b11111111011000011010100101111101;
   assign mem[7852] = 32'b00000000010100101111100010000000;
   assign mem[7853] = 32'b00000010110000011111111110011100;
   assign mem[7854] = 32'b00000101101101001110111010011000;
   assign mem[7855] = 32'b11111011100111100010011000001000;
   assign mem[7856] = 32'b11110110001001011100000001010000;
   assign mem[7857] = 32'b11111101000101101010011010111100;
   assign mem[7858] = 32'b00000001110000111110000100100000;
   assign mem[7859] = 32'b00000100011001110100111100111000;
   assign mem[7860] = 32'b11111011110110101111011100100000;
   assign mem[7861] = 32'b11111101011100101011101110000000;
   assign mem[7862] = 32'b11111110001100100101101001000110;
   assign mem[7863] = 32'b11111111011001110101101000100011;
   assign mem[7864] = 32'b00001000101101011001100111010000;
   assign mem[7865] = 32'b00001010011010111100000001100000;
   assign mem[7866] = 32'b11111111100010001101111101101100;
   assign mem[7867] = 32'b00000001111111000001101101111010;
   assign mem[7868] = 32'b11111001010110000001000111011000;
   assign mem[7869] = 32'b11111110001101100111111101111100;
   assign mem[7870] = 32'b11101111010110111100101100100000;
   assign mem[7871] = 32'b11101111101010111010111100000000;
   assign mem[7872] = 32'b00000100011101000010101010000000;
   assign mem[7873] = 32'b00001001110111011101000101110000;
   assign mem[7874] = 32'b11111101010111001111111010001000;
   assign mem[7875] = 32'b00000000001001000000101100100011;
   assign mem[7876] = 32'b11111011010110000101111011001000;
   assign mem[7877] = 32'b00000000101001000011011001110100;
   assign mem[7878] = 32'b00000101101110110010010001100000;
   assign mem[7879] = 32'b00000101010100111101100101000000;
   assign mem[7880] = 32'b11111000010000010000011101101000;
   assign mem[7881] = 32'b00000101101100011111101011100000;
   assign mem[7882] = 32'b11111011101010110001011000010000;
   assign mem[7883] = 32'b11111110001101110000111010110010;
   assign mem[7884] = 32'b11111111000110100100011110001001;
   assign mem[7885] = 32'b00000000000110000100011111000110;
   assign mem[7886] = 32'b11111111110010110011000101111011;
   assign mem[7887] = 32'b00001001000111110101101000000000;
   assign mem[7888] = 32'b11111110100101011111110111100010;
   assign mem[7889] = 32'b00000000100000010011001000101101;
   assign mem[7890] = 32'b11110101101110101010010001000000;
   assign mem[7891] = 32'b11111011100110110010111001000000;
   assign mem[7892] = 32'b00000011110100011010010010111100;
   assign mem[7893] = 32'b00000011001000111111101000100100;
   assign mem[7894] = 32'b00000001010101110001101001001010;
   assign mem[7895] = 32'b00000010010110100111000011010100;
   assign mem[7896] = 32'b00000000111010101000000111101110;
   assign mem[7897] = 32'b11110111000110101010110110100000;
   assign mem[7898] = 32'b00000101001111100110010110101000;
   assign mem[7899] = 32'b00000110111101110110101100110000;
   assign mem[7900] = 32'b00000011011101101001001111110100;
   assign mem[7901] = 32'b00000010110100011110110111100100;
   assign mem[7902] = 32'b11111110100000010010101111000010;
   assign mem[7903] = 32'b00000001100111000110111101010100;
   assign mem[7904] = 32'b00000001100111010000110100011000;
   assign mem[7905] = 32'b11111100101100100101011000000100;
   assign mem[7906] = 32'b00000101010000111011110100101000;
   assign mem[7907] = 32'b11111000001101110000010110001000;
   assign mem[7908] = 32'b00000001011001100110000101101110;
   assign mem[7909] = 32'b11111111101011011011111001000101;
   assign mem[7910] = 32'b11111100011100111111000001011100;
   assign mem[7911] = 32'b00000011101100111110000111011100;
   assign mem[7912] = 32'b11110010111101011000001101010000;
   assign mem[7913] = 32'b00000101000011110010101101011000;
   assign mem[7914] = 32'b11111011001000101111111100111000;
   assign mem[7915] = 32'b00000001110111110111101001110100;
   assign mem[7916] = 32'b11111100101010111100111010001100;
   assign mem[7917] = 32'b11111010000001011101110100111000;
   assign mem[7918] = 32'b00001000100011100010110010110000;
   assign mem[7919] = 32'b11111111011000100011010100110011;
   assign mem[7920] = 32'b11111110000010000101100001011100;
   assign mem[7921] = 32'b00000000001011110111100011111010;
   assign mem[7922] = 32'b11110110010010100001000100110000;
   assign mem[7923] = 32'b00000000000110011000011110001001;
   assign mem[7924] = 32'b11111110101001011100100111000100;
   assign mem[7925] = 32'b00000100011110011010110101111000;
   assign mem[7926] = 32'b11110101110100000011001100000000;
   assign mem[7927] = 32'b11111001100011110000010001010000;
   assign mem[7928] = 32'b00001011011010010000011100010000;
   assign mem[7929] = 32'b00000000101010111011000010111011;
   assign mem[7930] = 32'b00000001000111001010010111010010;
   assign mem[7931] = 32'b00000111100001100101000011111000;
   assign mem[7932] = 32'b11111101101011000101011110000100;
   assign mem[7933] = 32'b11110000100010110001100111100000;
   assign mem[7934] = 32'b11111100100111011010110001000000;
   assign mem[7935] = 32'b00000101010011100110011100100000;
   assign mem[7936] = 32'b00000000100101000001001011011001;
   assign mem[7937] = 32'b00001100011101010001101000110000;
   assign mem[7938] = 32'b11110111100110011000100100010000;
   assign mem[7939] = 32'b11111011111011100111000011101000;
   assign mem[7940] = 32'b00001001010001101011000001110000;
   assign mem[7941] = 32'b11111010000100101100101110010000;
   assign mem[7942] = 32'b11110101100000000011011001010000;
   assign mem[7943] = 32'b11101110011001110100101101100000;
   assign mem[7944] = 32'b00000100111001100011111011011000;
   assign mem[7945] = 32'b00000001011000100101001100101110;
   assign mem[7946] = 32'b00000001011001000010100110101000;
   assign mem[7947] = 32'b00000110011011110101100101001000;
   assign mem[7948] = 32'b00000110110011100100100100110000;
   assign mem[7949] = 32'b11111111011000110101101001110000;
   assign mem[7950] = 32'b11110001011110111010100000110000;
   assign mem[7951] = 32'b00001001111010111101000110100000;
   assign mem[7952] = 32'b00000100000010101001100011010000;
   assign mem[7953] = 32'b00000000000000100111110100111010;
   assign mem[7954] = 32'b11111000000101111000101101000000;
   assign mem[7955] = 32'b11111010001001100100000010110000;
   assign mem[7956] = 32'b00001010001101110111001001100000;
   assign mem[7957] = 32'b00000111000101000111010011011000;
   assign mem[7958] = 32'b11111010100000100111001101011000;
   assign mem[7959] = 32'b11111100010001110111000001110100;
   assign mem[7960] = 32'b11110100001000100110001001100000;
   assign mem[7961] = 32'b11101011100011110100010111000000;
   assign mem[7962] = 32'b11111101111010010011111001000100;
   assign mem[7963] = 32'b00000000000111111000101100001001;
   assign mem[7964] = 32'b00001001110011100111011000110000;
   assign mem[7965] = 32'b00000100000111101100100011101000;
   assign mem[7966] = 32'b00000000101010101110010101010101;
   assign mem[7967] = 32'b11110001111011111101101010110000;
   assign mem[7968] = 32'b00000001101011111101111111011100;
   assign mem[7969] = 32'b00000110001111100110000100001000;
   assign mem[7970] = 32'b11101100110001101000001000000000;
   assign mem[7971] = 32'b00000000100101100011010001010101;
   assign mem[7972] = 32'b00000111111001000100010001111000;
   assign mem[7973] = 32'b00000010101111000100111000101100;
   assign mem[7974] = 32'b00000110001010111000011100101000;
   assign mem[7975] = 32'b00000101110101110001100100111000;
   assign mem[7976] = 32'b00000101010111101010010011100000;
   assign mem[7977] = 32'b00001000100110001100110000010000;
   assign mem[7978] = 32'b11111000111011110110100001000000;
   assign mem[7979] = 32'b11110111111100100011000101110000;
   assign mem[7980] = 32'b00000100100001111001111010110000;
   assign mem[7981] = 32'b00001000001100111011001110010000;
   assign mem[7982] = 32'b11111110101001101111111101001100;
   assign mem[7983] = 32'b11111001011011110011101111000000;
   assign mem[7984] = 32'b11111011000111010111001101111000;
   assign mem[7985] = 32'b00000101110001011100000101100000;
   assign mem[7986] = 32'b11111111111111111111010111011011;
   assign mem[7987] = 32'b00000010000101100000011111101000;
   assign mem[7988] = 32'b11111111110010111101100001010010;
   assign mem[7989] = 32'b11110111010000110000000110000000;
   assign mem[7990] = 32'b00000010001000001101111010011000;
   assign mem[7991] = 32'b11101111001010100100011011000000;
   assign mem[7992] = 32'b11110110101010010110000111110000;
   assign mem[7993] = 32'b11111110010111000100010000110100;
   assign mem[7994] = 32'b00000010000100001011001110001000;
   assign mem[7995] = 32'b00000011100101001010110101011000;
   assign mem[7996] = 32'b11111111011001010001110000001110;
   assign mem[7997] = 32'b00000010011001010000011101100000;
   assign mem[7998] = 32'b11111010111101000011011001011000;
   assign mem[7999] = 32'b00000111010001110000001100011000;
   assign mem[8000] = 32'b00000000010100101001100100100111;
   assign mem[8001] = 32'b11111110110011011000100101100110;
   assign mem[8002] = 32'b00000000110100100010011011110001;
   assign mem[8003] = 32'b00000010010000100010011100110000;
   assign mem[8004] = 32'b11111100001001001101100101100000;
   assign mem[8005] = 32'b11111101111001111001010001001000;
   assign mem[8006] = 32'b00000000101000111100010010101010;
   assign mem[8007] = 32'b11111111010001000110001001010110;
   assign mem[8008] = 32'b00000000100101011110111111111100;
   assign mem[8009] = 32'b11111100101100110010010001010100;
   assign mem[8010] = 32'b00000101001111001101100010100000;
   assign mem[8011] = 32'b00000011110001010001000011111000;
   assign mem[8012] = 32'b00000000011101110100100001110100;
   assign mem[8013] = 32'b00000010100111000110100111011100;
   assign mem[8014] = 32'b11111100111110111000101110001000;
   assign mem[8015] = 32'b00000000100100011001100011100000;
   assign mem[8016] = 32'b00000110011110101011001001001000;
   assign mem[8017] = 32'b00000011000101100011001000111100;
   assign mem[8018] = 32'b11111010100110000011100010110000;
   assign mem[8019] = 32'b11111000001101010011111000100000;
   assign mem[8020] = 32'b11111110100100110111010001010100;
   assign mem[8021] = 32'b11111011001000110110011101110000;
   assign mem[8022] = 32'b11111101010001101110101011101100;
   assign mem[8023] = 32'b11111100110011111010001010001000;
   assign mem[8024] = 32'b00000111001011110100001110110000;
   assign mem[8025] = 32'b00000010111101011000000011000100;
   assign mem[8026] = 32'b00000010100011100010110111011100;
   assign mem[8027] = 32'b11111011011110011101100110000000;
   assign mem[8028] = 32'b11111100001000010000000011010100;
   assign mem[8029] = 32'b00000010100100100000101110101100;
   assign mem[8030] = 32'b00000100011111101001110100111000;
   assign mem[8031] = 32'b00000010100100011000111110110000;
   assign mem[8032] = 32'b11111011100011100000101010001000;
   assign mem[8033] = 32'b00001010101010101000001111100000;
   assign mem[8034] = 32'b11111111101111111001100001111010;
   assign mem[8035] = 32'b11111110101011010010010000001010;
   assign mem[8036] = 32'b11111111010001000011010010100101;
   assign mem[8037] = 32'b00010010010011110110110101100000;
   assign mem[8038] = 32'b11100110000111100001000000000000;
   assign mem[8039] = 32'b11111011000010010000000010110000;
   assign mem[8040] = 32'b11111010100101000011100100111000;
   assign mem[8041] = 32'b11100100000011111100011110100000;
   assign mem[8042] = 32'b00000110111101111110001011111000;
   assign mem[8043] = 32'b11111101011011000101110101101100;
   assign mem[8044] = 32'b00000101001000111011000000111000;
   assign mem[8045] = 32'b00000100001010111000110011100000;
   assign mem[8046] = 32'b11111110011111101110110100010000;
   assign mem[8047] = 32'b11111100011100111110101000100000;
   assign mem[8048] = 32'b00000000001101111110111101101010;
   assign mem[8049] = 32'b11111011011001001011110111111000;
   assign mem[8050] = 32'b11110110011110101100000001110000;
   assign mem[8051] = 32'b00000011001110000011000101001000;
   assign mem[8052] = 32'b00000100011000000100010110001000;
   assign mem[8053] = 32'b11111100011110111111001101011000;
   assign mem[8054] = 32'b00000011101100110100111000001100;
   assign mem[8055] = 32'b00000100110000011010110001101000;
   assign mem[8056] = 32'b00000001100011101100011011111110;
   assign mem[8057] = 32'b11110101000111010011010000010000;
   assign mem[8058] = 32'b00000001110100011001111011000000;
   assign mem[8059] = 32'b11111110000100010000111101100000;
   assign mem[8060] = 32'b11111100111011111100110011110000;
   assign mem[8061] = 32'b11110110111001110010101101100000;
   assign mem[8062] = 32'b11110011101111011000101101000000;
   assign mem[8063] = 32'b11111101110100100000011000100000;
   assign mem[8064] = 32'b00000110100011001011001010011000;
   assign mem[8065] = 32'b00000011110101011100001000000100;
   assign mem[8066] = 32'b00000001011110000110110100011110;
   assign mem[8067] = 32'b11110000010100011010100000100000;
   assign mem[8068] = 32'b00000101000000000001001011011000;
   assign mem[8069] = 32'b00000110011010000101011110010000;
   assign mem[8070] = 32'b11111010101000000001100100000000;
   assign mem[8071] = 32'b00000000010000101110110010001101;
   assign mem[8072] = 32'b00000101110100101000111000100000;
   assign mem[8073] = 32'b00000111110011000100110110100000;
   assign mem[8074] = 32'b11110011011011110100101001100000;
   assign mem[8075] = 32'b11110111111001000101110100000000;
   assign mem[8076] = 32'b11111000010111011101011111001000;
   assign mem[8077] = 32'b00000110011000101000010001001000;
   assign mem[8078] = 32'b11101111110000111111111111100000;
   assign mem[8079] = 32'b00000000110001110001110001000011;
   assign mem[8080] = 32'b00001001001001100100011101000000;
   assign mem[8081] = 32'b00000101010110010000101101011000;
   assign mem[8082] = 32'b11111001001001000000000000111000;
   assign mem[8083] = 32'b11111001001001011101010110111000;
   assign mem[8084] = 32'b00000100101000010110000111000000;
   assign mem[8085] = 32'b11111011110011011111000010100000;
   assign mem[8086] = 32'b11110111010010100010010000100000;
   assign mem[8087] = 32'b11111110010000000101111101110100;
   assign mem[8088] = 32'b00000101010110000000101100010000;
   assign mem[8089] = 32'b11111110110111100111011000000010;
   assign mem[8090] = 32'b11111111110100001011111101111000;
   assign mem[8091] = 32'b11110110111101001101000101000000;
   assign mem[8092] = 32'b00000010100100111011101100101000;
   assign mem[8093] = 32'b00000100111010101001101111010000;
   assign mem[8094] = 32'b11111101111110011110101001110000;
   assign mem[8095] = 32'b00000001100100101001100000001010;
   assign mem[8096] = 32'b00000001000101010010011100111100;
   assign mem[8097] = 32'b00000010100011011011111110101100;
   assign mem[8098] = 32'b11111001101110100010110001111000;
   assign mem[8099] = 32'b11111101101000110001010101110000;
   assign mem[8100] = 32'b00000001110100101100101011011110;
   assign mem[8101] = 32'b11110101111111011001001100010000;
   assign mem[8102] = 32'b00001000000011110010100110010000;
   assign mem[8103] = 32'b00001000000110110110110110010000;
   assign mem[8104] = 32'b11111100100100001011111100100100;
   assign mem[8105] = 32'b00000100010101111100101011110000;
   assign mem[8106] = 32'b11101011100000001001010010100000;
   assign mem[8107] = 32'b11111101100010101011111101000000;
   assign mem[8108] = 32'b11101011000100001101001101100000;
   assign mem[8109] = 32'b00000110100001001111111101111000;
   assign mem[8110] = 32'b00001011011001111010011000010000;
   assign mem[8111] = 32'b00000100110111100011110110000000;
   assign mem[8112] = 32'b11111101101010000101110100111000;
   assign mem[8113] = 32'b11101111001001001010000101000000;
   assign mem[8114] = 32'b00000000100000111111001101011101;
   assign mem[8115] = 32'b00001000001101111111011100110000;
   assign mem[8116] = 32'b11111110010011010110010101110100;
   assign mem[8117] = 32'b11111011110000011110000000110000;
   assign mem[8118] = 32'b00000001010100111100111110110000;
   assign mem[8119] = 32'b11110100000011001101101001010000;
   assign mem[8120] = 32'b11111110100110111000001101101110;
   assign mem[8121] = 32'b11111010110000110100011001110000;
   assign mem[8122] = 32'b11111001101010111101111101111000;
   assign mem[8123] = 32'b00000001000100110011011111010000;
   assign mem[8124] = 32'b00000100011010001100111101011000;
   assign mem[8125] = 32'b00000010101101011100011000110100;
   assign mem[8126] = 32'b00000010101100100000110010011100;
   assign mem[8127] = 32'b11101101111100111011110101000000;
   assign mem[8128] = 32'b00000001100011110111101010110010;
   assign mem[8129] = 32'b00001000011111110001001001000000;
   assign mem[8130] = 32'b11101101101000010000101011100000;
   assign mem[8131] = 32'b00001001011010111011100100110000;
   assign mem[8132] = 32'b00000101101110001101101010011000;
   assign mem[8133] = 32'b11110011011101010111111100000000;
   assign mem[8134] = 32'b11111100010000100110101110011000;
   assign mem[8135] = 32'b00000011010010011100011000000100;
   assign mem[8136] = 32'b11110111000011000101011110100000;
   assign mem[8137] = 32'b11111000101111100101111111000000;
   assign mem[8138] = 32'b00001101000010010101110000000000;
   assign mem[8139] = 32'b11111100111100100111010111100000;
   assign mem[8140] = 32'b11111101110000100001100111001100;
   assign mem[8141] = 32'b00000010011000100110011010101000;
   assign mem[8142] = 32'b11111101110111000001111011000100;
   assign mem[8143] = 32'b11111011100101110101001000110000;
   assign mem[8144] = 32'b00000011000011001101010000011000;
   assign mem[8145] = 32'b00000000100111000001111101111010;
   assign mem[8146] = 32'b11110111100110111111001101110000;
   assign mem[8147] = 32'b11111111101000000011000011011011;
   assign mem[8148] = 32'b11111101111101110101110011010100;
   assign mem[8149] = 32'b00000100001011110010101001101000;
   assign mem[8150] = 32'b00000011010011101111111111110000;
   assign mem[8151] = 32'b11111111011110101001001010101111;
   assign mem[8152] = 32'b00000011000111100011110101111100;
   assign mem[8153] = 32'b00000000001010111110001011011000;
   assign mem[8154] = 32'b00000010111010000111000110111100;
   assign mem[8155] = 32'b11111111010010001001101101001110;
   assign mem[8156] = 32'b00000011000101110000111111111100;
   assign mem[8157] = 32'b11111110110000000001011100111000;
   assign mem[8158] = 32'b11111011110001100101000111010000;
   assign mem[8159] = 32'b11111101010110001100110011001100;
   assign mem[8160] = 32'b00000010101000010010001011000100;
   assign mem[8161] = 32'b00000001001110011110001111011100;
   assign mem[8162] = 32'b11111000100011001111110000010000;
   assign mem[8163] = 32'b11111101101011110001110011100000;
   assign mem[8164] = 32'b00000000111111111110000100000010;
   assign mem[8165] = 32'b00000011111111110100101000101100;
   assign mem[8166] = 32'b00000001110111100100110011101100;
   assign mem[8167] = 32'b00000010100111100101101111110000;
   assign mem[8168] = 32'b00000010100000101011110110001100;
   assign mem[8169] = 32'b11111100001111111110000101010000;
   assign mem[8170] = 32'b11111001000001111100010010110000;
   assign mem[8171] = 32'b00000101010010001111000110000000;
   assign mem[8172] = 32'b00000000011000101110100110000011;
   assign mem[8173] = 32'b00000111000000110000110000101000;
   assign mem[8174] = 32'b11110011100010110001111000000000;
   assign mem[8175] = 32'b00000010110010101110110010010100;
   assign mem[8176] = 32'b00000101101101100100011111010000;
   assign mem[8177] = 32'b00000110001000110000001110011000;
   assign mem[8178] = 32'b11111011011000010110010000011000;
   assign mem[8179] = 32'b11111010001111111000001110000000;
   assign mem[8180] = 32'b11111100011010010111000100011000;
   assign mem[8181] = 32'b11111010111010101000010011011000;
   assign mem[8182] = 32'b00000000111001000111110100011001;
   assign mem[8183] = 32'b11111101010111111010000111000100;
   assign mem[8184] = 32'b11111011101110111110100110101000;
   assign mem[8185] = 32'b11111011001010000010011110000000;
   assign mem[8186] = 32'b00000010011001111000010011110100;
   assign mem[8187] = 32'b11111101001000111000001101101000;
   assign mem[8188] = 32'b00000101011111011111001000110000;
   assign mem[8189] = 32'b00000111011011000011010101100000;
   assign mem[8190] = 32'b11111011011001111001111110101000;
   assign mem[8191] = 32'b00000100100001010101101110000000;
   assign mem[8192] = 32'b00000000111110010001011100100100;
   assign mem[8193] = 32'b00000000110011110100111100111001;
   assign mem[8194] = 32'b11111000101000111001111111000000;
   assign mem[8195] = 32'b11111111001110100111001101100111;
   assign mem[8196] = 32'b11111010101111100110100100100000;
   assign mem[8197] = 32'b00000110101111001010110111100000;
   assign mem[8198] = 32'b11111101101111001000001111110000;
   assign mem[8199] = 32'b11111000100111101110001010111000;
   assign mem[8200] = 32'b11111001001000100010010010100000;
   assign mem[8201] = 32'b11110100011011101110110111100000;
   assign mem[8202] = 32'b11110111101111011010010000010000;
   assign mem[8203] = 32'b00000011011110111000000001111000;
   assign mem[8204] = 32'b00001000101010100010010010000000;
   assign mem[8205] = 32'b11111110011010111011111011100110;
   assign mem[8206] = 32'b11111100011010001001001000000000;
   assign mem[8207] = 32'b00000000010100101010000000111110;
   assign mem[8208] = 32'b11111110000010111100110010100000;
   assign mem[8209] = 32'b00000111111010110100010111101000;
   assign mem[8210] = 32'b11110100001100000001000001110000;
   assign mem[8211] = 32'b11101111100111010110001101100000;
   assign mem[8212] = 32'b00000000101101011101001010110011;
   assign mem[8213] = 32'b00000011001110010011110001001100;
   assign mem[8214] = 32'b00000111010010001010011111010000;
   assign mem[8215] = 32'b00000010111111010101101010111000;
   assign mem[8216] = 32'b00000100010011111001101000011000;
   assign mem[8217] = 32'b11110101000110101101000011000000;
   assign mem[8218] = 32'b11111111101111011101111111000001;
   assign mem[8219] = 32'b00000001010000111110010011101100;
   assign mem[8220] = 32'b11111101100110100110001101010000;
   assign mem[8221] = 32'b00000001101110111001010000010110;
   assign mem[8222] = 32'b11111010000101000100010100101000;
   assign mem[8223] = 32'b00000110010101100010101011101000;
   assign mem[8224] = 32'b11111110111111111110101000100000;
   assign mem[8225] = 32'b00000011001100000001000001100100;
   assign mem[8226] = 32'b11111110100000101010110000010010;
   assign mem[8227] = 32'b00000010011001110100010111010100;
   assign mem[8228] = 32'b11111100010001111010100110001000;
   assign mem[8229] = 32'b11111110001000100111100010100010;
   assign mem[8230] = 32'b00000100000111001100110111000000;
   assign mem[8231] = 32'b00000001101000000010110000001010;
   assign mem[8232] = 32'b11110101110111010011011111000000;
   assign mem[8233] = 32'b11111001101000010001011010110000;
   assign mem[8234] = 32'b00000011010010100100101011000000;
   assign mem[8235] = 32'b11111110111000111001001000100000;
   assign mem[8236] = 32'b00000000111000010011101110001111;
   assign mem[8237] = 32'b00000101100111001111110101011000;
   assign mem[8238] = 32'b11110011111101100110010000100000;
   assign mem[8239] = 32'b00000100001110010101001011110000;
   assign mem[8240] = 32'b00000110111001101000110101111000;
   assign mem[8241] = 32'b00001010010110011010011111100000;
   assign mem[8242] = 32'b11111011101100100000010100110000;
   assign mem[8243] = 32'b00000100001000000010011111011000;
   assign mem[8244] = 32'b11111010110111010100100010111000;
   assign mem[8245] = 32'b11111110010100111110101111100000;
   assign mem[8246] = 32'b11111001101101000101111100011000;
   assign mem[8247] = 32'b11111001101010110101100001101000;
   assign mem[8248] = 32'b11111011010011001100101010111000;
   assign mem[8249] = 32'b00000000010010010001110101111100;
   assign mem[8250] = 32'b11111101101101100010101000100100;
   assign mem[8251] = 32'b11111010010000010100000110101000;
   assign mem[8252] = 32'b11111100011000101001101000011100;
   assign mem[8253] = 32'b11111100101010100111000010110000;
   assign mem[8254] = 32'b00000010100100111011110011000100;
   assign mem[8255] = 32'b00000000011001011111110111001001;
   assign mem[8256] = 32'b11110001101010001001000110110000;
   assign mem[8257] = 32'b11111100111101100110000001000100;
   assign mem[8258] = 32'b00000111100010010111011100100000;
   assign mem[8259] = 32'b00000100100110001101101010110000;
   assign mem[8260] = 32'b11111010011001110100100001110000;
   assign mem[8261] = 32'b11111000010001010010001010110000;
   assign mem[8262] = 32'b00001100111010011001000010010000;
   assign mem[8263] = 32'b11111010010111011110011000111000;
   assign mem[8264] = 32'b11111011001111011110010001101000;
   assign mem[8265] = 32'b00001000010111010101011011000000;
   assign mem[8266] = 32'b00001001000110110101101011010000;
   assign mem[8267] = 32'b00000011011101110010001100110100;
   assign mem[8268] = 32'b11111001101110001111000110011000;
   assign mem[8269] = 32'b11110110111000110111011011000000;
   assign mem[8270] = 32'b11111011010100000101001000110000;
   assign mem[8271] = 32'b00000010100010011101100111111000;
   assign mem[8272] = 32'b00000100010100100110001001101000;
   assign mem[8273] = 32'b11110110011110111010101010000000;
   assign mem[8274] = 32'b11111100011100011100010111101100;
   assign mem[8275] = 32'b00000001000011011100011101011100;
   assign mem[8276] = 32'b00000001010111110000111111010000;
   assign mem[8277] = 32'b11111010110101100001001011011000;
   assign mem[8278] = 32'b00001101000000100010001101010000;
   assign mem[8279] = 32'b11111010010010110011100000101000;
   assign mem[8280] = 32'b11110100011001001010101100010000;
   assign mem[8281] = 32'b00000000101001100011110101100000;
   assign mem[8282] = 32'b00001000011011100011110010000000;
   assign mem[8283] = 32'b00001000010000101110000000000000;
   assign mem[8284] = 32'b11110111100010110000101011010000;
   assign mem[8285] = 32'b11111110010110010001100011010000;
   assign mem[8286] = 32'b00001010110000111010110011010000;
   assign mem[8287] = 32'b00000011011110010011000000001000;
   assign mem[8288] = 32'b11110110001100100010100101000000;
   assign mem[8289] = 32'b11111110010100101111001100001100;
   assign mem[8290] = 32'b00000001100100001001101110110100;
   assign mem[8291] = 32'b00000100111001000010111100111000;
   assign mem[8292] = 32'b00000000111110111011101100010010;
   assign mem[8293] = 32'b00000011110010101010000110101100;
   assign mem[8294] = 32'b11110110111100011110011000010000;
   assign mem[8295] = 32'b00000001010010100011110111101010;
   assign mem[8296] = 32'b00001000011000100110001010000000;
   assign mem[8297] = 32'b00000000111101000111011001000010;
   assign mem[8298] = 32'b11110110101100000111010111010000;
   assign mem[8299] = 32'b11110111010011000100000110000000;
   assign mem[8300] = 32'b11101010011111111100011100000000;
   assign mem[8301] = 32'b00000110110010100100011011110000;
   assign mem[8302] = 32'b11111000100110101001010011111000;
   assign mem[8303] = 32'b00000010001111011101011111010100;
   assign mem[8304] = 32'b11110101101000111100001001110000;
   assign mem[8305] = 32'b00000110111110010010100010000000;
   assign mem[8306] = 32'b00000000011010000010010001011110;
   assign mem[8307] = 32'b00000110111110101010111000001000;
   assign mem[8308] = 32'b11111111111110110101000100111110;
   assign mem[8309] = 32'b11110111000110111011010010000000;
   assign mem[8310] = 32'b11101110111001111010000110000000;
   assign mem[8311] = 32'b00000011011110010001000000011100;
   assign mem[8312] = 32'b00000000010100011001010111111010;
   assign mem[8313] = 32'b11111000101010100011011111010000;
   assign mem[8314] = 32'b11110001111100001001000111010000;
   assign mem[8315] = 32'b00000001110001000100010111101100;
   assign mem[8316] = 32'b11111111100100001010101001011001;
   assign mem[8317] = 32'b00001000111010010111010110100000;
   assign mem[8318] = 32'b00000010110101001011110001111100;
   assign mem[8319] = 32'b11111001101001111111011011011000;
   assign mem[8320] = 32'b00000000011001010110111001110101;
   assign mem[8321] = 32'b11110110011011111011010111110000;
   assign mem[8322] = 32'b11111111111100100100101101010111;
   assign mem[8323] = 32'b00001011111111000000111000000000;
   assign mem[8324] = 32'b11111101110001011001101001110100;
   assign mem[8325] = 32'b11111010111100010001111001001000;
   assign mem[8326] = 32'b00000111000010011101011100010000;
   assign mem[8327] = 32'b00000100101111110110011010100000;
   assign mem[8328] = 32'b00001000000101101111010100010000;
   assign mem[8329] = 32'b11110101101001010011100101010000;
   assign mem[8330] = 32'b00000011000010011111000010011000;
   assign mem[8331] = 32'b00000100010011111110110001001000;
   assign mem[8332] = 32'b00000010010111000010110100010000;
   assign mem[8333] = 32'b00000010000010111000011001110000;
   assign mem[8334] = 32'b11110100110110100111001101110000;
   assign mem[8335] = 32'b00001000001101110111101100100000;
   assign mem[8336] = 32'b00000111100101001111101001010000;
   assign mem[8337] = 32'b11110110100110001000011010000000;
   assign mem[8338] = 32'b11101100100101011110011110000000;
   assign mem[8339] = 32'b00000101101011001000101100100000;
   assign mem[8340] = 32'b11111110001101111101101110001110;
   assign mem[8341] = 32'b11111111000010011111011011011011;
   assign mem[8342] = 32'b11110111101001000011110011010000;
   assign mem[8343] = 32'b00000100100101110100001110011000;
   assign mem[8344] = 32'b11110110100010101101111001000000;
   assign mem[8345] = 32'b00000101010000101000000010110000;
   assign mem[8346] = 32'b00000101101100011111011100101000;
   assign mem[8347] = 32'b11111110110101011011111010101110;
   assign mem[8348] = 32'b00000000101010011011101011100111;
   assign mem[8349] = 32'b11111110011110101111001101010100;
   assign mem[8350] = 32'b00000010010011111001100101110100;
   assign mem[8351] = 32'b11110111111000001000101000110000;
   assign mem[8352] = 32'b11110101110111010111010111010000;
   assign mem[8353] = 32'b00000111000101111101110100111000;
   assign mem[8354] = 32'b11110000101111001110100010100000;
   assign mem[8355] = 32'b00000110100111110111110110100000;
   assign mem[8356] = 32'b11111010011111110101100000101000;
   assign mem[8357] = 32'b00000010011111010001000101001100;
   assign mem[8358] = 32'b00000000000010110100111011000011;
   assign mem[8359] = 32'b00000010001101000111110101001100;
   assign mem[8360] = 32'b11111110111010111000000100101010;
   assign mem[8361] = 32'b11110011100010011000100101000000;
   assign mem[8362] = 32'b11111110011101101111101001000010;
   assign mem[8363] = 32'b11111010011011011111000110101000;
   assign mem[8364] = 32'b11110010101010110000011110100000;
   assign mem[8365] = 32'b00000100111001100011111100001000;
   assign mem[8366] = 32'b11111001001001100100110100111000;
   assign mem[8367] = 32'b00000001100001010011010001000100;
   assign mem[8368] = 32'b11111100111011001001100011110000;
   assign mem[8369] = 32'b00000101010000111000110101000000;
   assign mem[8370] = 32'b11111100000111110101001110001100;
   assign mem[8371] = 32'b00000100000001100011011011001000;
   assign mem[8372] = 32'b00000110010110000110000110010000;
   assign mem[8373] = 32'b00000001001101100100101000110010;
   assign mem[8374] = 32'b11111111010111001100010001110100;
   assign mem[8375] = 32'b11100111110100100011010010100000;
   assign mem[8376] = 32'b11111010001010010000011000011000;
   assign mem[8377] = 32'b00000100000011111000001110001000;
   assign mem[8378] = 32'b00000010110111011100010000000100;
   assign mem[8379] = 32'b11111001101011111010111000100000;
   assign mem[8380] = 32'b00000001010001000010000001100100;
   assign mem[8381] = 32'b00000000001101110000101100101011;
   assign mem[8382] = 32'b11111111000111111011111000110011;
   assign mem[8383] = 32'b11110110110001000010110110000000;
   assign mem[8384] = 32'b11111001101001101111001000011000;
   assign mem[8385] = 32'b00000100110100001100100010001000;
   assign mem[8386] = 32'b11111110100011001000110110010110;
   assign mem[8387] = 32'b00000011100001001011000111000100;
   assign mem[8388] = 32'b11111110011010111110111000001010;
   assign mem[8389] = 32'b00000111101111111010000000001000;
   assign mem[8390] = 32'b11110101000001001110100110100000;
   assign mem[8391] = 32'b11111111101100011100110101101001;
   assign mem[8392] = 32'b00000101010100010111010101101000;
   assign mem[8393] = 32'b00000110101010111110011001110000;
   assign mem[8394] = 32'b11111110010111010001100101000010;
   assign mem[8395] = 32'b11101101000010001110100000100000;
   assign mem[8396] = 32'b11111010110100010011111011100000;
   assign mem[8397] = 32'b00000100101111111000000010010000;
   assign mem[8398] = 32'b00000001011000010011010000100000;
   assign mem[8399] = 32'b11111111000110000011001011010101;
   assign mem[8400] = 32'b11110011101101000011101111100000;
   assign mem[8401] = 32'b11111110001010011101011111011100;
   assign mem[8402] = 32'b00000101100001000101101011000000;
   assign mem[8403] = 32'b11110111011111100001010011110000;
   assign mem[8404] = 32'b11110101111100110010100111000000;
   assign mem[8405] = 32'b00001000000000001000101001100000;
   assign mem[8406] = 32'b00000111111101111100101000110000;
   assign mem[8407] = 32'b11110001101110011001110111010000;
   assign mem[8408] = 32'b11110011001011100011000101110000;
   assign mem[8409] = 32'b00000100101001011010100001111000;
   assign mem[8410] = 32'b00000010011111110001001101101100;
   assign mem[8411] = 32'b11111011100101001000000010000000;
   assign mem[8412] = 32'b00001000000001111001100110010000;
   assign mem[8413] = 32'b11101010101000010000101110000000;
   assign mem[8414] = 32'b00000010111100110011010100010100;
   assign mem[8415] = 32'b00000111101111000111000111001000;
   assign mem[8416] = 32'b11110101011101100110111110110000;
   assign mem[8417] = 32'b00001001111000011000000101000000;
   assign mem[8418] = 32'b11110001110110101001000111100000;
   assign mem[8419] = 32'b11111010100010011111000111100000;
   assign mem[8420] = 32'b11101011101111111101111011000000;
   assign mem[8421] = 32'b11111010001000111111100000110000;
   assign mem[8422] = 32'b11111001101011001101111001010000;
   assign mem[8423] = 32'b00000010000101001001011000111100;
   assign mem[8424] = 32'b00000011011010100111101110010100;
   assign mem[8425] = 32'b00000001011110001100000000101010;
   assign mem[8426] = 32'b00000101110110101010100110001000;
   assign mem[8427] = 32'b00000110011110111011011000110000;
   assign mem[8428] = 32'b00000101110110100001001010111000;
   assign mem[8429] = 32'b00000010101001100100110101011000;
   assign mem[8430] = 32'b00000101110000011001001110101000;
   assign mem[8431] = 32'b11111111110111010000100000001101;
   assign mem[8432] = 32'b11111100000100100010010100111000;
   assign mem[8433] = 32'b00000000010001111011001011110011;
   assign mem[8434] = 32'b11111011001111011100011111001000;
   assign mem[8435] = 32'b11111110010111101111001011001000;
   assign mem[8436] = 32'b00000000110001001000001110100000;
   assign mem[8437] = 32'b00000100001001101101101011011000;
   assign mem[8438] = 32'b00000000000110100010111010110100;
   assign mem[8439] = 32'b00000000000110110011101110110000;
   assign mem[8440] = 32'b11110100111111110001001111110000;
   assign mem[8441] = 32'b11110011011101111011111101110000;
   assign mem[8442] = 32'b00000101100011011100001110111000;
   assign mem[8443] = 32'b00000011010110100000110000001100;
   assign mem[8444] = 32'b00000110001100100011010101101000;
   assign mem[8445] = 32'b00000001001100101010101110010010;
   assign mem[8446] = 32'b00000100010010000111011110101000;
   assign mem[8447] = 32'b00001011001110011111110100010000;
   assign mem[8448] = 32'b00000010000101100001011010100000;
   assign mem[8449] = 32'b11110000010000000100111111100000;
   assign mem[8450] = 32'b11110000100111101000111100100000;
   assign mem[8451] = 32'b11110111001001000010100000000000;
   assign mem[8452] = 32'b11111101111010110100100011011100;
   assign mem[8453] = 32'b00000011101010011100111100001000;
   assign mem[8454] = 32'b11111000001010110010100101110000;
   assign mem[8455] = 32'b00000100001101000011111101000000;
   assign mem[8456] = 32'b00001000010010001101101010100000;
   assign mem[8457] = 32'b11111110111101010000001111100110;
   assign mem[8458] = 32'b11111111010011101011110011010011;
   assign mem[8459] = 32'b11111001000000001100000111000000;
   assign mem[8460] = 32'b11111001101001111011010110101000;
   assign mem[8461] = 32'b11110111000010110111101000110000;
   assign mem[8462] = 32'b11111011111100111010001010010000;
   assign mem[8463] = 32'b00000100001111111011110110110000;
   assign mem[8464] = 32'b00000010010001101001110000001000;
   assign mem[8465] = 32'b11111011110011010110110011111000;
   assign mem[8466] = 32'b00000010010010101001101101000100;
   assign mem[8467] = 32'b11111110001011010111000000010100;
   assign mem[8468] = 32'b00000010000001101000111011111000;
   assign mem[8469] = 32'b00000011110010100011011111010000;
   assign mem[8470] = 32'b00000010111111111000011000101100;
   assign mem[8471] = 32'b11111101111110101111100110011100;
   assign mem[8472] = 32'b00000101011110000011100110000000;
   assign mem[8473] = 32'b11111101110011110010010110001100;
   assign mem[8474] = 32'b00000010111110110000101101000100;
   assign mem[8475] = 32'b11110110111101000101001110000000;
   assign mem[8476] = 32'b11111001001111100111111100001000;
   assign mem[8477] = 32'b00000011110010000000111101001000;
   assign mem[8478] = 32'b00000000010010011111110011110010;
   assign mem[8479] = 32'b11111010000011100100111101010000;
   assign mem[8480] = 32'b11110011111110101000110101000000;
   assign mem[8481] = 32'b11110111110111100101110010010000;
   assign mem[8482] = 32'b11111101011001111011111000011100;
   assign mem[8483] = 32'b00000110100011001101011000010000;
   assign mem[8484] = 32'b00001011100101011110010000000000;
   assign mem[8485] = 32'b11110111111001011100100000100000;
   assign mem[8486] = 32'b11110101111111000010110011100000;
   assign mem[8487] = 32'b11111111010001111010111110000011;
   assign mem[8488] = 32'b00001000010010010110101011110000;
   assign mem[8489] = 32'b00000111100110111011001010111000;
   assign mem[8490] = 32'b11110110111011101010111001110000;
   assign mem[8491] = 32'b11111011100110100110100110100000;
   assign mem[8492] = 32'b11111101110001110110000111011100;
   assign mem[8493] = 32'b00000010001101000111100010001100;
   assign mem[8494] = 32'b00000111110101011111011111111000;
   assign mem[8495] = 32'b00000000100111101010111011101011;
   assign mem[8496] = 32'b11111111000110111010011110011101;
   assign mem[8497] = 32'b11111100110111100100100011001000;
   assign mem[8498] = 32'b11111101001000101110000101111100;
   assign mem[8499] = 32'b00000100101110001110001111100000;
   assign mem[8500] = 32'b11111101001001001110010011010100;
   assign mem[8501] = 32'b11110110011100110001011101010000;
   assign mem[8502] = 32'b11111001101110001000100001010000;
   assign mem[8503] = 32'b00000100011010001011111010001000;
   assign mem[8504] = 32'b11110001000000101101010100010000;
   assign mem[8505] = 32'b00000111100101000011010000011000;
   assign mem[8506] = 32'b00001000010011111010000001000000;
   assign mem[8507] = 32'b11111011110100100100110000001000;
   assign mem[8508] = 32'b11111111000000110110010111011000;
   assign mem[8509] = 32'b00000000011001001001000011000101;
   assign mem[8510] = 32'b11111110110110000101010011011000;
   assign mem[8511] = 32'b11101000100110100010100111100000;
   assign mem[8512] = 32'b11111100101000001000001110010000;
   assign mem[8513] = 32'b00000110100011101101111001101000;
   assign mem[8514] = 32'b11111010101101001001011111010000;
   assign mem[8515] = 32'b11111011110010100100011110110000;
   assign mem[8516] = 32'b00000110101010101100010100110000;
   assign mem[8517] = 32'b11111111110001100011001010000111;
   assign mem[8518] = 32'b00000000000010000001011011110011;
   assign mem[8519] = 32'b00000010010000011110001001101000;
   assign mem[8520] = 32'b00000010001001010101010000011100;
   assign mem[8521] = 32'b00000001111100111000110000010010;
   assign mem[8522] = 32'b00000100010000011100111011110000;
   assign mem[8523] = 32'b11110101011100011010100001100000;
   assign mem[8524] = 32'b00000010101010101101010011011100;
   assign mem[8525] = 32'b11111101110000110011100101001100;
   assign mem[8526] = 32'b11111011011011000010101100110000;
   assign mem[8527] = 32'b00000101011000110010110010111000;
   assign mem[8528] = 32'b11110110001011011110101100000000;
   assign mem[8529] = 32'b00000000010000000010011100001101;
   assign mem[8530] = 32'b11111000000110101011001001111000;
   assign mem[8531] = 32'b11111010001011101001011000011000;
   assign mem[8532] = 32'b11111101110110100111010000101000;
   assign mem[8533] = 32'b00000010000101001000000001101000;
   assign mem[8534] = 32'b11111010001001100100111000010000;
   assign mem[8535] = 32'b00000001000010010010011100111110;
   assign mem[8536] = 32'b00000100101010111110001111100000;
   assign mem[8537] = 32'b11111110110100000110111011110100;
   assign mem[8538] = 32'b00000111001100000010111010100000;
   assign mem[8539] = 32'b00000110010101000011110000100000;
   assign mem[8540] = 32'b11111100001110010010100101101000;
   assign mem[8541] = 32'b11111110101011111100010011011100;
   assign mem[8542] = 32'b00000010011001101101101000101100;
   assign mem[8543] = 32'b00001001011010110011110100110000;
   assign mem[8544] = 32'b11111101101100001101001010111100;
   assign mem[8545] = 32'b11110000010000010000110100100000;
   assign mem[8546] = 32'b11111001100110010001110111000000;
   assign mem[8547] = 32'b00000010011011100100111011000000;
   assign mem[8548] = 32'b00000101010110110111010000010000;
   assign mem[8549] = 32'b00000001010011100101110011001010;
   assign mem[8550] = 32'b00000100111101101100100001101000;
   assign mem[8551] = 32'b00000000100101110111011100111111;
   assign mem[8552] = 32'b11111100010011011111011111111100;
   assign mem[8553] = 32'b00000001001010101110011100010110;
   assign mem[8554] = 32'b00001001000011100111100000100000;
   assign mem[8555] = 32'b00000000000000111011100100101010;
   assign mem[8556] = 32'b11110111011010111110000100100000;
   assign mem[8557] = 32'b00000101110001110100101010001000;
   assign mem[8558] = 32'b11111111010010100000001111111000;
   assign mem[8559] = 32'b00000000100110110100100101110110;
   assign mem[8560] = 32'b00001010010011100110100000000000;
   assign mem[8561] = 32'b11111111110110011100100010101011;
   assign mem[8562] = 32'b00000010011000011001110100000100;
   assign mem[8563] = 32'b11111110001110111001010111110010;
   assign mem[8564] = 32'b00000011011011110000000111100000;
   assign mem[8565] = 32'b11111110111101101111101011110110;
   assign mem[8566] = 32'b11111100010011100000011110001100;
   assign mem[8567] = 32'b00000101110000010010011111110000;
   assign mem[8568] = 32'b11111011111011110001010111001000;
   assign mem[8569] = 32'b00000000000111001111110110001010;
   assign mem[8570] = 32'b11111000010111100000000100000000;
   assign mem[8571] = 32'b00000000001010011111011100010011;
   assign mem[8572] = 32'b00000001000110100101011011000010;
   assign mem[8573] = 32'b00000001011110010111101101010000;
   assign mem[8574] = 32'b11111100110010111101001101110100;
   assign mem[8575] = 32'b11111110000110100010011100101100;
   assign mem[8576] = 32'b11111001100001111100010011111000;
   assign mem[8577] = 32'b00000010111111100011000101100000;
   assign mem[8578] = 32'b11111111000100101110011100100110;
   assign mem[8579] = 32'b00000011100010000001100111011000;
   assign mem[8580] = 32'b00000010000110110011001001000000;
   assign mem[8581] = 32'b00000010111110101000000001110100;
   assign mem[8582] = 32'b11111101111100000010001100001100;
   assign mem[8583] = 32'b11111011000011010101111001011000;
   assign mem[8584] = 32'b00000100101010101010000110010000;
   assign mem[8585] = 32'b11110101000111111010001011000000;
   assign mem[8586] = 32'b11111011111011011000101110011000;
   assign mem[8587] = 32'b00000001101111000101010111010000;
   assign mem[8588] = 32'b00000000011010001011010110100110;
   assign mem[8589] = 32'b11111110101000011011001011100110;
   assign mem[8590] = 32'b11111110100011011011111110110100;
   assign mem[8591] = 32'b11111111011001000111000101110110;
   assign mem[8592] = 32'b00001001000000011011000000000000;
   assign mem[8593] = 32'b11101100011101100001101010100000;
   assign mem[8594] = 32'b00000011001000001100111000100000;
   assign mem[8595] = 32'b11111110110000100001000111110010;
   assign mem[8596] = 32'b00000010000111010001100001111100;
   assign mem[8597] = 32'b11111001111001001000101101010000;
   assign mem[8598] = 32'b00000111111011000000101101110000;
   assign mem[8599] = 32'b11111100101011000011011010001100;
   assign mem[8600] = 32'b11110100010010101110001001000000;
   assign mem[8601] = 32'b11101101001010100001100010100000;
   assign mem[8602] = 32'b11111100010100110011110110000000;
   assign mem[8603] = 32'b00000100000100011101000110000000;
   assign mem[8604] = 32'b00000110000111100100101100110000;
   assign mem[8605] = 32'b11110110101001000011001010110000;
   assign mem[8606] = 32'b00000010111001000000000000001000;
   assign mem[8607] = 32'b11111100110101001110000010001100;
   assign mem[8608] = 32'b00000100011111101100010100001000;
   assign mem[8609] = 32'b00000011110000010111010100011100;
   assign mem[8610] = 32'b11110110100001010111100111000000;
   assign mem[8611] = 32'b11111010001101000100111101101000;
   assign mem[8612] = 32'b00001001010011101111001000110000;
   assign mem[8613] = 32'b11111100110101000100011011100000;
   assign mem[8614] = 32'b11110110010010011110011010100000;
   assign mem[8615] = 32'b00000110100111010111000000110000;
   assign mem[8616] = 32'b00001110110001011110111101100000;
   assign mem[8617] = 32'b11111111011100010001110010001000;
   assign mem[8618] = 32'b11110101110110111000101001000000;
   assign mem[8619] = 32'b11111011101011110000000110101000;
   assign mem[8620] = 32'b00000101100011001111000100110000;
   assign mem[8621] = 32'b00000110011100001001100111001000;
   assign mem[8622] = 32'b00000000011010011011001010111000;
   assign mem[8623] = 32'b11111101100001110100000100110100;
   assign mem[8624] = 32'b00000000111111011010011000000010;
   assign mem[8625] = 32'b11111111110111010110010110011011;
   assign mem[8626] = 32'b11110001011110110000101110010000;
   assign mem[8627] = 32'b00000100010110100000011010101000;
   assign mem[8628] = 32'b11111110010010101011101100000010;
   assign mem[8629] = 32'b11111110010001110010110100110100;
   assign mem[8630] = 32'b00000011001010101011101010111100;
   assign mem[8631] = 32'b11101110000110110011010000100000;
   assign mem[8632] = 32'b11110110110010001100010001100000;
   assign mem[8633] = 32'b00000010111010011001101010111100;
   assign mem[8634] = 32'b00000001001111110000101100011110;
   assign mem[8635] = 32'b11111110000011011101111101001010;
   assign mem[8636] = 32'b00000000101000010000001110101010;
   assign mem[8637] = 32'b00001011100110010011100110100000;
   assign mem[8638] = 32'b00000100001011101000110100010000;
   assign mem[8639] = 32'b11111010011110100111000010111000;
   assign mem[8640] = 32'b11110010001010101010010000110000;
   assign mem[8641] = 32'b00000111111010010010110000011000;
   assign mem[8642] = 32'b00000000100010001100100110001011;
   assign mem[8643] = 32'b00001010100010000010001110000000;
   assign mem[8644] = 32'b11111111011110100101100010101110;
   assign mem[8645] = 32'b11101000010011000001010101000000;
   assign mem[8646] = 32'b11111011000111101010111011011000;
   assign mem[8647] = 32'b11111110100100110111101111010100;
   assign mem[8648] = 32'b00000101001010101001001111011000;
   assign mem[8649] = 32'b00000010001100010110001001001100;
   assign mem[8650] = 32'b11111101111111011011110101110000;
   assign mem[8651] = 32'b00000011101000001101010000101100;
   assign mem[8652] = 32'b00000100111111001000111111001000;
   assign mem[8653] = 32'b11110101001100001100100010110000;
   assign mem[8654] = 32'b11111111010000001101100101001100;
   assign mem[8655] = 32'b11111000111000010100000001101000;
   assign mem[8656] = 32'b11111110110010100111010001100100;
   assign mem[8657] = 32'b00000111100100101111001000111000;
   assign mem[8658] = 32'b00000101000000110010000111000000;
   assign mem[8659] = 32'b11110111110000011110000101010000;
   assign mem[8660] = 32'b11110110110001001100000100110000;
   assign mem[8661] = 32'b11111110110011000000110001000010;
   assign mem[8662] = 32'b11111100000110001001110111101100;
   assign mem[8663] = 32'b00000101100111111111010110110000;
   assign mem[8664] = 32'b00000010001110001111011011001100;
   assign mem[8665] = 32'b00000001110110110111110100010100;
   assign mem[8666] = 32'b11111111111100010011000100101001;
   assign mem[8667] = 32'b00000110001111010111010001001000;
   assign mem[8668] = 32'b11111111111010001101000001100000;
   assign mem[8669] = 32'b11111001011010011110111111100000;
   assign mem[8670] = 32'b00000101010001001100011000110000;
   assign mem[8671] = 32'b00000101010100101010110111111000;
   assign mem[8672] = 32'b00000100001111011011001111111000;
   assign mem[8673] = 32'b11111001001101100001100010001000;
   assign mem[8674] = 32'b11111001010000000000100001110000;
   assign mem[8675] = 32'b11110101111101100011010001000000;
   assign mem[8676] = 32'b11111100111001110111100011010100;
   assign mem[8677] = 32'b00000000010110110110100101010000;
   assign mem[8678] = 32'b11111100000011011110000000001000;
   assign mem[8679] = 32'b00000011111011010100000100001000;
   assign mem[8680] = 32'b11110111111110001011100100100000;
   assign mem[8681] = 32'b11101110001110111100000010100000;
   assign mem[8682] = 32'b00000100000100010000001100001000;
   assign mem[8683] = 32'b00000111000001100100011011111000;
   assign mem[8684] = 32'b11111101111010000110111110011000;
   assign mem[8685] = 32'b00000110010010000010010011000000;
   assign mem[8686] = 32'b00001010011001000110010001000000;
   assign mem[8687] = 32'b11101111011001110100111101100000;
   assign mem[8688] = 32'b00000001010001111010000101010000;
   assign mem[8689] = 32'b11110111000110000110001100100000;
   assign mem[8690] = 32'b11111000001011000111111010110000;
   assign mem[8691] = 32'b11111011110110000010111111011000;
   assign mem[8692] = 32'b11111001001001000110010100010000;
   assign mem[8693] = 32'b00000001111011111110001011100000;
   assign mem[8694] = 32'b11111100011011111110111011111000;
   assign mem[8695] = 32'b00000100100001101110110000001000;
   assign mem[8696] = 32'b00000110111010100110101000111000;
   assign mem[8697] = 32'b11111010100000110101100011001000;
   assign mem[8698] = 32'b00000001010010101110110000010000;
   assign mem[8699] = 32'b11111111010001110010111101111101;
   assign mem[8700] = 32'b11111101100010001100101110000000;
   assign mem[8701] = 32'b11111110110101000110010100110110;
   assign mem[8702] = 32'b11111011101010000110100001110000;
   assign mem[8703] = 32'b00000101000100001010000001111000;
   assign mem[8704] = 32'b00000100010111010010000010000000;
   assign mem[8705] = 32'b11110101011000001110010110000000;
   assign mem[8706] = 32'b11110101011101100001010010100000;
   assign mem[8707] = 32'b00001001100010110001000000000000;
   assign mem[8708] = 32'b00001001101011001000011011110000;
   assign mem[8709] = 32'b00000100100100001000100111111000;
   assign mem[8710] = 32'b11111001111110010110010000111000;
   assign mem[8711] = 32'b11110111101111010111010000000000;
   assign mem[8712] = 32'b00000011100000101111111011001100;
   assign mem[8713] = 32'b11111110111010010011011011011010;
   assign mem[8714] = 32'b11110110011101100100010001000000;
   assign mem[8715] = 32'b11111100111111010101111100100000;
   assign mem[8716] = 32'b11111110010001110111111000101000;
   assign mem[8717] = 32'b11111110100000101111101011010110;
   assign mem[8718] = 32'b00000111110000110011011010110000;
   assign mem[8719] = 32'b00000010100010101000111100101100;
   assign mem[8720] = 32'b00000000110000001100011101100001;
   assign mem[8721] = 32'b00000100011101101010000011000000;
   assign mem[8722] = 32'b11110111110000000101100111100000;
   assign mem[8723] = 32'b00000010101100011111101101101100;
   assign mem[8724] = 32'b11111111101011100011101111010011;
   assign mem[8725] = 32'b00000100011111011100001011010000;
   assign mem[8726] = 32'b11111101111100000111001100011100;
   assign mem[8727] = 32'b00000011110101011111011100010100;
   assign mem[8728] = 32'b11111111011001100000011001011100;
   assign mem[8729] = 32'b11111111111000100001000011011110;
   assign mem[8730] = 32'b11111100010111101111001010010100;
   assign mem[8731] = 32'b11111010111001010011001100100000;
   assign mem[8732] = 32'b11111001111000011110100000000000;
   assign mem[8733] = 32'b00000111010010111110000000001000;
   assign mem[8734] = 32'b00000001110011000011111010010110;
   assign mem[8735] = 32'b11111111100110011110110010000101;
   assign mem[8736] = 32'b11110111100011000110100110100000;
   assign mem[8737] = 32'b11111011110101110101111000010000;
   assign mem[8738] = 32'b00000100000111011101101100100000;
   assign mem[8739] = 32'b00001010110111010011001111000000;
   assign mem[8740] = 32'b00001100100110011110100010100000;
   assign mem[8741] = 32'b11111111110000000001001110110100;
   assign mem[8742] = 32'b11101101100011101111100100100000;
   assign mem[8743] = 32'b11111110110001110101100011100010;
   assign mem[8744] = 32'b11101111101110011010101100100000;
   assign mem[8745] = 32'b00000110100010000100010100000000;
   assign mem[8746] = 32'b11111010011110111010110001111000;
   assign mem[8747] = 32'b00010000011001100000111000000000;
   assign mem[8748] = 32'b11110001000110011001101011100000;
   assign mem[8749] = 32'b11111101111010000001100011001000;
   assign mem[8750] = 32'b00000001011110110100000001011000;
   assign mem[8751] = 32'b00000010100000001010111110000100;
   assign mem[8752] = 32'b00000000100101010111011110010111;
   assign mem[8753] = 32'b11111111000000000000001111011011;
   assign mem[8754] = 32'b11111110101011010010101010100100;
   assign mem[8755] = 32'b11111000011111000000100001101000;
   assign mem[8756] = 32'b11111100011100101111001111011000;
   assign mem[8757] = 32'b11111110100011111100110011001110;
   assign mem[8758] = 32'b11111100011101000010010110100000;
   assign mem[8759] = 32'b00000001111010101001111001010000;
   assign mem[8760] = 32'b11111001000000010100010010100000;
   assign mem[8761] = 32'b00000101101110010101101101010000;
   assign mem[8762] = 32'b11111011111001001111000101000000;
   assign mem[8763] = 32'b00000010011010011100010101000100;
   assign mem[8764] = 32'b00001010100101101111001000110000;
   assign mem[8765] = 32'b11111001000000000000101110011000;
   assign mem[8766] = 32'b11110110000110100000001010100000;
   assign mem[8767] = 32'b00001010000100011100010000110000;
   assign mem[8768] = 32'b11111000000100010001000110001000;
   assign mem[8769] = 32'b11111110101100011000101010011010;
   assign mem[8770] = 32'b00000000001000101001000001011011;
   assign mem[8771] = 32'b11111110111101111011011110001010;
   assign mem[8772] = 32'b00000010011100110111101100101000;
   assign mem[8773] = 32'b00000100010110111110011111011000;
   assign mem[8774] = 32'b11111011000111000000011001010000;
   assign mem[8775] = 32'b00000100100000110010000110001000;
   assign mem[8776] = 32'b00000110010111011100001111111000;
   assign mem[8777] = 32'b11111000000001101111001110011000;
   assign mem[8778] = 32'b00000000101111000101000110000011;
   assign mem[8779] = 32'b11111111101101000111110111010110;
   assign mem[8780] = 32'b11111111110100000100010100001111;
   assign mem[8781] = 32'b11111011010111011000110100111000;
   assign mem[8782] = 32'b00000001001000000011001010001000;
   assign mem[8783] = 32'b11111110101001011100101011010100;
   assign mem[8784] = 32'b11111111111101001011111110001010;
   assign mem[8785] = 32'b00000010100100111100001100110000;
   assign mem[8786] = 32'b11110111101111110000011100110000;
   assign mem[8787] = 32'b00001000001001011000000110000000;
   assign mem[8788] = 32'b11111001010101000010111010101000;
   assign mem[8789] = 32'b11111001111101010100100000010000;
   assign mem[8790] = 32'b00000100001011110001000101110000;
   assign mem[8791] = 32'b00000000000110110010111111000000;
   assign mem[8792] = 32'b00000000111101011101100100100000;
   assign mem[8793] = 32'b11111100001111100100000001110000;
   assign mem[8794] = 32'b00000010010011110010011100111100;
   assign mem[8795] = 32'b00000010101100111101011011110100;
   assign mem[8796] = 32'b00000010100111101111010111111100;
   assign mem[8797] = 32'b11111101100011101010111010010100;
   assign mem[8798] = 32'b00000001111101100110110110110100;
   assign mem[8799] = 32'b11111100011111010100110011010100;
   assign mem[8800] = 32'b11110110111001001010101100010000;
   assign mem[8801] = 32'b00000111000011000001111000101000;
   assign mem[8802] = 32'b11111110001011110011000001111110;
   assign mem[8803] = 32'b00000111000111101001010001101000;
   assign mem[8804] = 32'b00000010100101110000000001100000;
   assign mem[8805] = 32'b11111101101010110111110000100000;
   assign mem[8806] = 32'b00000000111100000010010100001001;
   assign mem[8807] = 32'b00000000111110001101100011001100;
   assign mem[8808] = 32'b00000001000100010011110000010110;
   assign mem[8809] = 32'b00001001001010101111111001100000;
   assign mem[8810] = 32'b11111111111000101010010100011111;
   assign mem[8811] = 32'b00000000101011111011110101110100;
   assign mem[8812] = 32'b11111101101110111011111000011000;
   assign mem[8813] = 32'b11110100110110110110000011100000;
   assign mem[8814] = 32'b00000000110110001000000111001010;
   assign mem[8815] = 32'b11110100011000110110110010110000;
   assign mem[8816] = 32'b00000011010010111000100111011000;
   assign mem[8817] = 32'b11111111101111011000111001101011;
   assign mem[8818] = 32'b00000101100100111110010001100000;
   assign mem[8819] = 32'b00000010000100100101100111000100;
   assign mem[8820] = 32'b11111111011010111100011111011010;
   assign mem[8821] = 32'b11111011010110010110001010011000;
   assign mem[8822] = 32'b00000000100000111011001001001101;
   assign mem[8823] = 32'b00000000110011011001010111101110;
   assign mem[8824] = 32'b00000001000100001101111111010110;
   assign mem[8825] = 32'b11110000100100001100000001100000;
   assign mem[8826] = 32'b11111011000001011011011011101000;
   assign mem[8827] = 32'b00000010010011001001111010011100;
   assign mem[8828] = 32'b00000100100111001000100011100000;
   assign mem[8829] = 32'b00000000101011011000100111101101;
   assign mem[8830] = 32'b00000000001111101111100001100001;
   assign mem[8831] = 32'b00000111100101111100010001001000;
   assign mem[8832] = 32'b00010000100001100110100001100000;
   assign mem[8833] = 32'b11101111001100110111111110000000;
   assign mem[8834] = 32'b00001111100111011001100001010000;
   assign mem[8835] = 32'b00000011111001100011101100110100;
   assign mem[8836] = 32'b11101111000010100010110100000000;
   assign mem[8837] = 32'b00000010110111010001011001001000;
   assign mem[8838] = 32'b11110011010100000000111101010000;
   assign mem[8839] = 32'b11111011101001100111010000010000;
   assign mem[8840] = 32'b11110110001101110011011000010000;
   assign mem[8841] = 32'b11110101001001101000111111010000;
   assign mem[8842] = 32'b11111100110011001011111100110100;
   assign mem[8843] = 32'b00000111100111000000100101011000;
   assign mem[8844] = 32'b11111111001101011010000011011011;
   assign mem[8845] = 32'b00000000111001011010001001110000;
   assign mem[8846] = 32'b00000101100111011000110000101000;
   assign mem[8847] = 32'b00000100001010011010100000100000;
   assign mem[8848] = 32'b11111100010011101111110010101000;
   assign mem[8849] = 32'b00000010110101011001101001101100;
   assign mem[8850] = 32'b11110010011110010101010001010000;
   assign mem[8851] = 32'b11110011011110110001000101000000;
   assign mem[8852] = 32'b00000000011110000001111110010011;
   assign mem[8853] = 32'b00000101100101001000000001111000;
   assign mem[8854] = 32'b11111100100101010010010001100000;
   assign mem[8855] = 32'b00000010100101101100111010100000;
   assign mem[8856] = 32'b00000101011000100010011110101000;
   assign mem[8857] = 32'b11111101001110100011101011101100;
   assign mem[8858] = 32'b11111111010001000010111011010001;
   assign mem[8859] = 32'b00000001101001111001101110010010;
   assign mem[8860] = 32'b11101110001000100111010010100000;
   assign mem[8861] = 32'b00000001100100000000111001100110;
   assign mem[8862] = 32'b11111111011011000011111100010011;
   assign mem[8863] = 32'b00000011111111011111110001100100;
   assign mem[8864] = 32'b00000001000001010011110010100110;
   assign mem[8865] = 32'b11111001110100100010000110010000;
   assign mem[8866] = 32'b11110111111111111001100100010000;
   assign mem[8867] = 32'b11111100000111011001111111111100;
   assign mem[8868] = 32'b00000011010110011000100001000000;
   assign mem[8869] = 32'b00000011000010000100101110000000;
   assign mem[8870] = 32'b11111110110000010100110001010110;
   assign mem[8871] = 32'b00000001000011110011111011011010;
   assign mem[8872] = 32'b00000100000010000000101010111000;
   assign mem[8873] = 32'b00000010110010001011110011101100;
   assign mem[8874] = 32'b11111010111111001101000100111000;
   assign mem[8875] = 32'b11111010000011011101100011110000;
   assign mem[8876] = 32'b11111101011110010010011100010000;
   assign mem[8877] = 32'b00000001010010011011010111100110;
   assign mem[8878] = 32'b11111110000111001111000010011010;
   assign mem[8879] = 32'b11111111110100100111110001010000;
   assign mem[8880] = 32'b11111011101000010110111101010000;
   assign mem[8881] = 32'b00000011110010101010110000011100;
   assign mem[8882] = 32'b11111110010001001010101110101000;
   assign mem[8883] = 32'b00000000100000111001101110110010;
   assign mem[8884] = 32'b00000010111000010101111010110100;
   assign mem[8885] = 32'b00000001010000010111100011100000;
   assign mem[8886] = 32'b11111011011000100010110011000000;
   assign mem[8887] = 32'b11111011000000101011001101110000;
   assign mem[8888] = 32'b11110010101101110110111100000000;
   assign mem[8889] = 32'b00001001111011110101110111110000;
   assign mem[8890] = 32'b00000111110100101010110110001000;
   assign mem[8891] = 32'b11110011110010001110000100100000;
   assign mem[8892] = 32'b11111001010001011010010011000000;
   assign mem[8893] = 32'b00000011000101101101010010001100;
   assign mem[8894] = 32'b11110110101101011010010100010000;
   assign mem[8895] = 32'b00000010001101100111010100000100;
   assign mem[8896] = 32'b11111111000011101111101111110101;
   assign mem[8897] = 32'b00000101001000010011011000111000;
   assign mem[8898] = 32'b00000011011010100101011000010000;
   assign mem[8899] = 32'b11111110100100010011010110101110;
   assign mem[8900] = 32'b11111010011011011010011100010000;
   assign mem[8901] = 32'b00000111110100100110011001010000;
   assign mem[8902] = 32'b00000100001111000111010110111000;
   assign mem[8903] = 32'b11111000001001000100001000100000;
   assign mem[8904] = 32'b00000000111101010010100101001111;
   assign mem[8905] = 32'b00000001101001101111010111110110;
   assign mem[8906] = 32'b00001000000110010010010101100000;
   assign mem[8907] = 32'b11111000001111010101001010010000;
   assign mem[8908] = 32'b11110001001100011110010111000000;
   assign mem[8909] = 32'b11111110101011000001011001111110;
   assign mem[8910] = 32'b11111011010001000111010100111000;
   assign mem[8911] = 32'b11111011011100001110101110010000;
   assign mem[8912] = 32'b11111100010010000100000110111100;
   assign mem[8913] = 32'b11111110000001001100011100001010;
   assign mem[8914] = 32'b00000010011010011000111011110000;
   assign mem[8915] = 32'b00000010111000100110110001001100;
   assign mem[8916] = 32'b00000101010101011111000110011000;
   assign mem[8917] = 32'b11111100010111000110110010001100;
   assign mem[8918] = 32'b00000011111110010010101001000000;
   assign mem[8919] = 32'b00000000001101010011111110001111;
   assign mem[8920] = 32'b11111110000110000110001011100010;
   assign mem[8921] = 32'b11111010110100100001010111000000;
   assign mem[8922] = 32'b00000000001110110010100011010011;
   assign mem[8923] = 32'b00000000001000001010110001101100;
   assign mem[8924] = 32'b11111010100011100100010110110000;
   assign mem[8925] = 32'b11111011101010110110110101000000;
   assign mem[8926] = 32'b00000100000010111011000110001000;
   assign mem[8927] = 32'b11110111111000111010110010010000;
   assign mem[8928] = 32'b00000110101011001100011100101000;
   assign mem[8929] = 32'b00000011001011000110001101001100;
   assign mem[8930] = 32'b11110110011110000001100101010000;
   assign mem[8931] = 32'b00000101011100110110011000100000;
   assign mem[8932] = 32'b00000011011010011111001101011100;
   assign mem[8933] = 32'b11110011111000110011000101000000;
   assign mem[8934] = 32'b00000101001111010000101100010000;
   assign mem[8935] = 32'b11110111111011101101111100010000;
   assign mem[8936] = 32'b00000101100011011001111100110000;
   assign mem[8937] = 32'b00000100100011011111011010000000;
   assign mem[8938] = 32'b00000110111010110101011000000000;
   assign mem[8939] = 32'b11111100100111101111100101000000;
   assign mem[8940] = 32'b00000111101111001101101100101000;
   assign mem[8941] = 32'b00000000111011010111010000100000;
   assign mem[8942] = 32'b00000101001011111010110010101000;
   assign mem[8943] = 32'b11101010011011100101100110100000;
   assign mem[8944] = 32'b00001011000000000010010000010000;
   assign mem[8945] = 32'b11111100001000001000110000101000;
   assign mem[8946] = 32'b11110111110110001111111010110000;
   assign mem[8947] = 32'b00000110011000111000011110000000;
   assign mem[8948] = 32'b11100110001001001100110001100000;
   assign mem[8949] = 32'b11111110000001110101100010011010;
   assign mem[8950] = 32'b00000000011001001101101000101110;
   assign mem[8951] = 32'b00000001101101101001001101111100;
   assign mem[8952] = 32'b00000110000111100111001001011000;
   assign mem[8953] = 32'b11110100000100110011011011100000;
   assign mem[8954] = 32'b00001010101111011010010101110000;
   assign mem[8955] = 32'b11111110010100000011000101111000;
   assign mem[8956] = 32'b11110010100010010011111011110000;
   assign mem[8957] = 32'b00000011010111001101101010000100;
   assign mem[8958] = 32'b11111011010001011010101100101000;
   assign mem[8959] = 32'b11111111011100011110011111100111;
   assign mem[8960] = 32'b11111111111000011111100111100010;
   assign mem[8961] = 32'b11111000010110011010100010100000;
   assign mem[8962] = 32'b00000110010111001001011100010000;
   assign mem[8963] = 32'b00001100011111010111010110000000;
   assign mem[8964] = 32'b00000000001010000010101111000111;
   assign mem[8965] = 32'b11111001010001110011100010101000;
   assign mem[8966] = 32'b00000011011111011000000010000100;
   assign mem[8967] = 32'b11111101101001100011011110001100;
   assign mem[8968] = 32'b00000111110001101101001111111000;
   assign mem[8969] = 32'b11101001011110100000000010000000;
   assign mem[8970] = 32'b11111011101010000100001011110000;
   assign mem[8971] = 32'b11111100000000111000001010110000;
   assign mem[8972] = 32'b11111011001111000111111111010000;
   assign mem[8973] = 32'b00000001010101011000011110101100;
   assign mem[8974] = 32'b11111110001000101111110111100110;
   assign mem[8975] = 32'b00000100000000010010111011100000;
   assign mem[8976] = 32'b00000011010010111001000110100100;
   assign mem[8977] = 32'b11111100101001001010111111000100;
   assign mem[8978] = 32'b11111011000110001011001001001000;
   assign mem[8979] = 32'b00000000011000000000111111111101;
   assign mem[8980] = 32'b00000001111111101100100111010010;
   assign mem[8981] = 32'b11111010000111100011101010110000;
   assign mem[8982] = 32'b11110101001010000100000101000000;
   assign mem[8983] = 32'b00000010001001010011000001010000;
   assign mem[8984] = 32'b11111000110011100101111101011000;
   assign mem[8985] = 32'b00000100100011000000010010011000;
   assign mem[8986] = 32'b00000011001001011000000000110100;
   assign mem[8987] = 32'b11111111010001100111100100011010;
   assign mem[8988] = 32'b00000010100111010011000110100000;
   assign mem[8989] = 32'b11110010111001101111011111000000;
   assign mem[8990] = 32'b00000011001101001001011000100000;
   assign mem[8991] = 32'b00000000100110110000101110001100;
   assign mem[8992] = 32'b11111011010000100110010110101000;
   assign mem[8993] = 32'b00000001001110111110011110100000;
   assign mem[8994] = 32'b00000001110011010000111100110010;
   assign mem[8995] = 32'b00001011100010110100111011010000;
   assign mem[8996] = 32'b11111000000001000010101101100000;
   assign mem[8997] = 32'b11111001010000010110001110101000;
   assign mem[8998] = 32'b11111101100110100001101000100100;
   assign mem[8999] = 32'b11111010001110111011111111011000;
   assign mem[9000] = 32'b11101011110011101100110010000000;
   assign mem[9001] = 32'b00000011001101011011011011110100;
   assign mem[9002] = 32'b11111101101011010111101101110000;
   assign mem[9003] = 32'b11111110110111010011110110000000;
   assign mem[9004] = 32'b00000000001011100001100110111011;
   assign mem[9005] = 32'b00000111011110101000000100111000;
   assign mem[9006] = 32'b00000011101001100110100010110100;
   assign mem[9007] = 32'b11111001101010000001111111111000;
   assign mem[9008] = 32'b00000010110111011101110011001000;
   assign mem[9009] = 32'b11111100111100011111111011101100;
   assign mem[9010] = 32'b00000110110000111001110001011000;
   assign mem[9011] = 32'b11111000100011101110001100110000;
   assign mem[9012] = 32'b00001000100001000100110100100000;
   assign mem[9013] = 32'b11111000100100111111110111111000;
   assign mem[9014] = 32'b00000010110101111001101010111000;
   assign mem[9015] = 32'b11101100111101110110000110100000;
   assign mem[9016] = 32'b11111111010001100010010011110010;
   assign mem[9017] = 32'b00000011101101110010001100000000;
   assign mem[9018] = 32'b00000101001100000110000000011000;
   assign mem[9019] = 32'b00000000011001011000011110001111;
   assign mem[9020] = 32'b11111101100111011101100011010100;
   assign mem[9021] = 32'b00000000110111000011100010110010;
   assign mem[9022] = 32'b00000000111101010010101001101011;
   assign mem[9023] = 32'b00000111010000010001000111011000;
   assign mem[9024] = 32'b00000010111100001000110001100100;
   assign mem[9025] = 32'b11111010011011101010100100000000;
   assign mem[9026] = 32'b11111011010011110110111000011000;
   assign mem[9027] = 32'b00000001100000101100010011100000;
   assign mem[9028] = 32'b00000100111000100110100011010000;
   assign mem[9029] = 32'b00000000101010101111111101101001;
   assign mem[9030] = 32'b00001000111101001110101101100000;
   assign mem[9031] = 32'b11110110001110101111110001010000;
   assign mem[9032] = 32'b00000110010001001110011101010000;
   assign mem[9033] = 32'b11111111011101011011001100001000;
   assign mem[9034] = 32'b00000111110001101000011001010000;
   assign mem[9035] = 32'b11100101101010001101011110000000;
   assign mem[9036] = 32'b11101100011101101100011101100000;
   assign mem[9037] = 32'b00000011111110111011011011110000;
   assign mem[9038] = 32'b00001001011011110010000111010000;
   assign mem[9039] = 32'b00000000000000001101111101001100;
   assign mem[9040] = 32'b11110010000000001000011100110000;
   assign mem[9041] = 32'b00000001110001100100110100110000;
   assign mem[9042] = 32'b00000001011100001101101111110100;
   assign mem[9043] = 32'b00000110010011100100010101001000;
   assign mem[9044] = 32'b11111000110010111001010111010000;
   assign mem[9045] = 32'b00000100000100101000111100001000;
   assign mem[9046] = 32'b00001000011100011011000000100000;
   assign mem[9047] = 32'b00000001110000100000010111100100;
   assign mem[9048] = 32'b11111100110111101001111001000100;
   assign mem[9049] = 32'b11111000011001010000000111110000;
   assign mem[9050] = 32'b00000000000101001100110011111000;
   assign mem[9051] = 32'b11111111010101111010010000100011;
   assign mem[9052] = 32'b00000000011010010000100111000110;
   assign mem[9053] = 32'b00000000101000111000111001101110;
   assign mem[9054] = 32'b11110010011111110100010000000000;
   assign mem[9055] = 32'b11110111111010001110111110110000;
   assign mem[9056] = 32'b11111001001011010101111001111000;
   assign mem[9057] = 32'b00000100100111010001010100101000;
   assign mem[9058] = 32'b00000100110111110111010100011000;
   assign mem[9059] = 32'b11111110101010110000111010111110;
   assign mem[9060] = 32'b00000001011011110101010101001010;
   assign mem[9061] = 32'b11110001110011111000110011010000;
   assign mem[9062] = 32'b00000100000110111010101100011000;
   assign mem[9063] = 32'b11110100100101110000100100110000;
   assign mem[9064] = 32'b00001011000010000100001101010000;
   assign mem[9065] = 32'b11110100010100010011111100010000;
   assign mem[9066] = 32'b00001001110110000111110111000000;
   assign mem[9067] = 32'b00000010011110110111100010111000;
   assign mem[9068] = 32'b00000011100111100110010011100000;
   assign mem[9069] = 32'b11110000100000000011010001110000;
   assign mem[9070] = 32'b00000101101010011110000101001000;
   assign mem[9071] = 32'b00000010011010111000101101110000;
   assign mem[9072] = 32'b11101111111111111111100111000000;
   assign mem[9073] = 32'b00000011010011000101011010110000;
   assign mem[9074] = 32'b00000001001100001110000110001100;
   assign mem[9075] = 32'b00000101100101110011111101101000;
   assign mem[9076] = 32'b00000100100001011101010110101000;
   assign mem[9077] = 32'b11111101010101110101111000101100;
   assign mem[9078] = 32'b00000010000100011100110110000100;
   assign mem[9079] = 32'b11110011100111010111100101010000;
   assign mem[9080] = 32'b11101111111100000010101011100000;
   assign mem[9081] = 32'b11111011010000010011010001100000;
   assign mem[9082] = 32'b00000100111011000001111000000000;
   assign mem[9083] = 32'b00000010111001101010110100111000;
   assign mem[9084] = 32'b00000101111100010010110101001000;
   assign mem[9085] = 32'b00000000101100010111110111000000;
   assign mem[9086] = 32'b11111111010011000111011111010110;
   assign mem[9087] = 32'b00000101110110110110001011110000;
   assign mem[9088] = 32'b11111111111111001101011000000100;
   assign mem[9089] = 32'b11101010001101011100011011000000;
   assign mem[9090] = 32'b11110110111000010011111011000000;
   assign mem[9091] = 32'b11111100100111101110111101000100;
   assign mem[9092] = 32'b00000000011101001100101110001110;
   assign mem[9093] = 32'b00000110110000000011101011100000;
   assign mem[9094] = 32'b00000010111101000001100111100100;
   assign mem[9095] = 32'b00000100100001010100001101010000;
   assign mem[9096] = 32'b00000010100001010001000011010100;
   assign mem[9097] = 32'b00000011011001110010000101000100;
   assign mem[9098] = 32'b00000010001111010111011101111100;
   assign mem[9099] = 32'b11110101101000011001011100110000;
   assign mem[9100] = 32'b11111010011110100111001100000000;
   assign mem[9101] = 32'b11110110100011010010100111000000;
   assign mem[9102] = 32'b00000010001111000111000000011000;
   assign mem[9103] = 32'b00001000011101001110111010000000;
   assign mem[9104] = 32'b00001001001010000000000110000000;
   assign mem[9105] = 32'b11110111101110101011101001000000;
   assign mem[9106] = 32'b11111010100010010110110001011000;
   assign mem[9107] = 32'b00000011000100010101010100010100;
   assign mem[9108] = 32'b00000010111100000100101100110100;
   assign mem[9109] = 32'b11111011000010011011110001100000;
   assign mem[9110] = 32'b00000111000101000001100011011000;
   assign mem[9111] = 32'b11110011000001100110111101010000;
   assign mem[9112] = 32'b00001000101000011001100100100000;
   assign mem[9113] = 32'b11101011101111010001000101000000;
   assign mem[9114] = 32'b11111010001100010101110001101000;
   assign mem[9115] = 32'b11110011111000110101100001110000;
   assign mem[9116] = 32'b11111111001111001001101000011000;
   assign mem[9117] = 32'b00000010110100000010011001110000;
   assign mem[9118] = 32'b00000100010011001000001010010000;
   assign mem[9119] = 32'b11110010001110011011110101100000;
   assign mem[9120] = 32'b11111100011010101101100011101100;
   assign mem[9121] = 32'b00000000000010001110011101101110;
   assign mem[9122] = 32'b00000111100100010011001001001000;
   assign mem[9123] = 32'b11110001110110011010000010110000;
   assign mem[9124] = 32'b00000100100100110001010100101000;
   assign mem[9125] = 32'b00000000111111010100011101110110;
   assign mem[9126] = 32'b11111001111011111100111010111000;
   assign mem[9127] = 32'b00000000100000010100110111111101;
   assign mem[9128] = 32'b00001000110001100011001111000000;
   assign mem[9129] = 32'b11111101011111110000011011001000;
   assign mem[9130] = 32'b00000111000011000100000110010000;
   assign mem[9131] = 32'b11111100101011100001101000011000;
   assign mem[9132] = 32'b11111001001001111001011000101000;
   assign mem[9133] = 32'b00000010001101110111110011111000;
   assign mem[9134] = 32'b11111101011100001100100101100000;
   assign mem[9135] = 32'b11111111101010000011001001101000;
   assign mem[9136] = 32'b00000101010011101100011001011000;
   assign mem[9137] = 32'b11111111100101011000001001010100;
   assign mem[9138] = 32'b00000001000001001011110111010100;
   assign mem[9139] = 32'b11111111001101111011000000111101;
   assign mem[9140] = 32'b11101011011111011101111010000000;
   assign mem[9141] = 32'b11110011001100010100101000010000;
   assign mem[9142] = 32'b11110110001000001101001110000000;
   assign mem[9143] = 32'b00000110110001111001010010000000;
   assign mem[9144] = 32'b00000000000000010000110110011001;
   assign mem[9145] = 32'b00000111011110011001010000101000;
   assign mem[9146] = 32'b00000100001110001111010100000000;
   assign mem[9147] = 32'b11111110001000101011010000011100;
   assign mem[9148] = 32'b00000011110000001001000011111000;
   assign mem[9149] = 32'b11111110001000011011110110000000;
   assign mem[9150] = 32'b00000010110110100011001110010100;
   assign mem[9151] = 32'b11100011010000110111010110000000;
   assign mem[9152] = 32'b11111111110000100000001100001110;
   assign mem[9153] = 32'b00000101001111000111011111011000;
   assign mem[9154] = 32'b00000000010010001001000101111000;
   assign mem[9155] = 32'b11111111001101111011010011111101;
   assign mem[9156] = 32'b00000100111001100011011000011000;
   assign mem[9157] = 32'b11111100000000000001011111010000;
   assign mem[9158] = 32'b00000110011100001101011101101000;
   assign mem[9159] = 32'b11111010010001110101010001010000;
   assign mem[9160] = 32'b00001001001010000110011011000000;
   assign mem[9161] = 32'b11111100101100110111001010100100;
   assign mem[9162] = 32'b11111111010011100000110110110101;
   assign mem[9163] = 32'b11101011001111101011010110000000;
   assign mem[9164] = 32'b00001101001111101010011001000000;
   assign mem[9165] = 32'b11110000011111000100000100000000;
   assign mem[9166] = 32'b11111100000110011010000111111000;
   assign mem[9167] = 32'b00001110101101101011010111010000;
   assign mem[9168] = 32'b11101111010110010011001101100000;
   assign mem[9169] = 32'b11111010001010001100111100110000;
   assign mem[9170] = 32'b11111011001010110101001101000000;
   assign mem[9171] = 32'b11110110000001111101010010110000;
   assign mem[9172] = 32'b00000111101010001010001111000000;
   assign mem[9173] = 32'b11111100001101010000011001111100;
   assign mem[9174] = 32'b00000001100111111001011111101110;
   assign mem[9175] = 32'b11111111110000101010111111100001;
   assign mem[9176] = 32'b00000101000001110111100010101000;
   assign mem[9177] = 32'b11111001110000101100110010010000;
   assign mem[9178] = 32'b00000101010010000110001110000000;
   assign mem[9179] = 32'b11111001101101110001001010111000;
   assign mem[9180] = 32'b00000011110100010100111000101100;
   assign mem[9181] = 32'b11111000110010001010100010011000;
   assign mem[9182] = 32'b00000111010010111001101010011000;
   assign mem[9183] = 32'b00000001100101101111101110011000;
   assign mem[9184] = 32'b00000000101011000100011110101110;
   assign mem[9185] = 32'b11101111011101010101101101100000;
   assign mem[9186] = 32'b11110101111101001010001111010000;
   assign mem[9187] = 32'b00000011101000001000100011111100;
   assign mem[9188] = 32'b00001000111000101101100000110000;
   assign mem[9189] = 32'b11111110100100010011011000000110;
   assign mem[9190] = 32'b00000010001110111011110111111000;
   assign mem[9191] = 32'b11111100110010110011101001011000;
   assign mem[9192] = 32'b11111010001101110001100001110000;
   assign mem[9193] = 32'b00000011001001110011101110001000;
   assign mem[9194] = 32'b00000111111111101010101001001000;
   assign mem[9195] = 32'b00000010111010011010001000001000;
   assign mem[9196] = 32'b11111110011101000000001111010100;
   assign mem[9197] = 32'b11111110101101110110010110000000;
   assign mem[9198] = 32'b11111110111010000100010100101100;
   assign mem[9199] = 32'b00000100100110001100010101110000;
   assign mem[9200] = 32'b00000100100101110100011000100000;
   assign mem[9201] = 32'b00000000111101101100001101011011;
   assign mem[9202] = 32'b11111111001100100100110101010000;
   assign mem[9203] = 32'b11111111101110010000111001000011;
   assign mem[9204] = 32'b00000101000110111111011011001000;
   assign mem[9205] = 32'b11111111001010110000011010011010;
   assign mem[9206] = 32'b11111010011111010110110110110000;
   assign mem[9207] = 32'b00000010000111101100101111101100;
   assign mem[9208] = 32'b11111000011100011010000110010000;
   assign mem[9209] = 32'b11111111100101011001101011010101;
   assign mem[9210] = 32'b11111100101011010100101101011100;
   assign mem[9211] = 32'b00000001010000111010000100011010;
   assign mem[9212] = 32'b00000000001010111111100011101011;
   assign mem[9213] = 32'b00000010011011101111001111011100;
   assign mem[9214] = 32'b00000010010110011101101110010000;
   assign mem[9215] = 32'b11111110011111010101000011100100;
   assign mem[9216] = 32'b11111010101100101110010001111000;
   assign mem[9217] = 32'b00000000000101011001011111001001;
   assign mem[9218] = 32'b11111101000001110110110001100100;
   assign mem[9219] = 32'b00000010110111001100010100011000;
   assign mem[9220] = 32'b11111111000100101100000101001101;
   assign mem[9221] = 32'b00000010000000011001010110111000;
   assign mem[9222] = 32'b00000000101110010110011111011100;
   assign mem[9223] = 32'b00000001100110001101101000110010;
   assign mem[9224] = 32'b00000000110000001101111110100000;
   assign mem[9225] = 32'b11111100001011111001101010101000;
   assign mem[9226] = 32'b11110101101000010011100110110000;
   assign mem[9227] = 32'b00000010000011111110001011100100;
   assign mem[9228] = 32'b11111110101000100101100101100000;
   assign mem[9229] = 32'b11111110111011100101001110110100;
   assign mem[9230] = 32'b11110111011101000001101100100000;
   assign mem[9231] = 32'b00000100101010011011000001100000;
   assign mem[9232] = 32'b00000111110100010011100000010000;
   assign mem[9233] = 32'b00000001100111101010111110001110;
   assign mem[9234] = 32'b11111010111100111010010001110000;
   assign mem[9235] = 32'b11110111101011001011110101100000;
   assign mem[9236] = 32'b11110010000111010100101001100000;
   assign mem[9237] = 32'b11111111011100111010000001000111;
   assign mem[9238] = 32'b00001000010100111100001001110000;
   assign mem[9239] = 32'b00000110111001000110110010001000;
   assign mem[9240] = 32'b11111101000100100001011110110000;
   assign mem[9241] = 32'b11111000101100000111101100101000;
   assign mem[9242] = 32'b00000010000010111001110000010100;
   assign mem[9243] = 32'b00001000001110110110100110110000;
   assign mem[9244] = 32'b00000010001111111001111000011100;
   assign mem[9245] = 32'b11101101011001000111011100100000;
   assign mem[9246] = 32'b00000000100110001001010110001000;
   assign mem[9247] = 32'b00001000001111101001110100100000;
   assign mem[9248] = 32'b00000100000110110010101111001000;
   assign mem[9249] = 32'b11110101010011111111000010010000;
   assign mem[9250] = 32'b11110111000010000111110100000000;
   assign mem[9251] = 32'b00000001100001000001010100000000;
   assign mem[9252] = 32'b00000011010101010000001011100000;
   assign mem[9253] = 32'b00000101100100111011100110010000;
   assign mem[9254] = 32'b11110101101111110000100011000000;
   assign mem[9255] = 32'b00000011001011110001010101010100;
   assign mem[9256] = 32'b00001010000010101110011001000000;
   assign mem[9257] = 32'b11111110110110001011001100011100;
   assign mem[9258] = 32'b11111011001100101000110100000000;
   assign mem[9259] = 32'b11110100000100001111110001110000;
   assign mem[9260] = 32'b00000010100011100111001000101000;
   assign mem[9261] = 32'b11111011111100001011001101010000;
   assign mem[9262] = 32'b00000010111110111111111000001100;
   assign mem[9263] = 32'b11110111011100111001010100010000;
   assign mem[9264] = 32'b00000101011000011010000111010000;
   assign mem[9265] = 32'b11111101111011110111110101100100;
   assign mem[9266] = 32'b11111000110101110101110111101000;
   assign mem[9267] = 32'b00000000001111011001001111001100;
   assign mem[9268] = 32'b11111100111111110101100010110100;
   assign mem[9269] = 32'b00000010000010001101101110001000;
   assign mem[9270] = 32'b00000001101100110101111100010000;
   assign mem[9271] = 32'b11111101110111110110001011100000;
   assign mem[9272] = 32'b11111111010100111011110001010001;
   assign mem[9273] = 32'b11110101110100011111001111000000;
   assign mem[9274] = 32'b00000101001100010001001101110000;
   assign mem[9275] = 32'b00000010100100011111100010111000;
   assign mem[9276] = 32'b11111000001011101010110001111000;
   assign mem[9277] = 32'b11111111111010011110111110000100;
   assign mem[9278] = 32'b00000001101011001010110001011010;
   assign mem[9279] = 32'b11111110111010010000000011000000;
   assign mem[9280] = 32'b11111110100111110100100011110100;
   assign mem[9281] = 32'b11110111111011110101011100000000;
   assign mem[9282] = 32'b11111111111111001011001010001101;
   assign mem[9283] = 32'b00000001010000000001111111111000;
   assign mem[9284] = 32'b11111110100110011110101111110010;
   assign mem[9285] = 32'b11101100010100111111001100100000;
   assign mem[9286] = 32'b11111100010111001111001010100000;
   assign mem[9287] = 32'b00000000000100010110000110100101;
   assign mem[9288] = 32'b00001011101101000111110011010000;
   assign mem[9289] = 32'b11111110110011111101101010001100;
   assign mem[9290] = 32'b00001001111100101010000100100000;
   assign mem[9291] = 32'b11111010100110110111111010001000;
   assign mem[9292] = 32'b11111100100110010000110100100100;
   assign mem[9293] = 32'b11110000010100111111001011100000;
   assign mem[9294] = 32'b00001000000101010000111001110000;
   assign mem[9295] = 32'b11110101110111101011101011110000;
   assign mem[9296] = 32'b11111110010011010110111010011100;
   assign mem[9297] = 32'b00000011011100000101001110110100;
   assign mem[9298] = 32'b11111110001011010101001001010110;
   assign mem[9299] = 32'b11111000011010101111100110011000;
   assign mem[9300] = 32'b11111110010010000101001101001000;
   assign mem[9301] = 32'b00000011001100110110110010101100;
   assign mem[9302] = 32'b00000111001000110100110011110000;
   assign mem[9303] = 32'b11110100101100000101011001100000;
   assign mem[9304] = 32'b00000111010100101010001000001000;
   assign mem[9305] = 32'b11111000100010100011001010011000;
   assign mem[9306] = 32'b00000010011001100001101100110100;
   assign mem[9307] = 32'b00000100001011111000000000100000;
   assign mem[9308] = 32'b00000001010111110100010010111010;
   assign mem[9309] = 32'b11111010010101000100100100100000;
   assign mem[9310] = 32'b00000010001011011111001000101100;
   assign mem[9311] = 32'b11111110011010011100100111000110;
   assign mem[9312] = 32'b00000000000111000001110010001001;
   assign mem[9313] = 32'b00000010110010001011100100110100;
   assign mem[9314] = 32'b00000000010110100010011011000010;
   assign mem[9315] = 32'b11101110000011011000100110000000;
   assign mem[9316] = 32'b11110101100010001100010001000000;
   assign mem[9317] = 32'b00000011100010100011010000010100;
   assign mem[9318] = 32'b00000011110000100101011101101000;
   assign mem[9319] = 32'b00000010000001010100011000000100;
   assign mem[9320] = 32'b11111000100111011111110010110000;
   assign mem[9321] = 32'b11110100101000010100010101100000;
   assign mem[9322] = 32'b11111010011011100110010011010000;
   assign mem[9323] = 32'b00000101001101010111000100001000;
   assign mem[9324] = 32'b11111000111000101010011100011000;
   assign mem[9325] = 32'b00000011010100000110001100000100;
   assign mem[9326] = 32'b00000101111010101100010001000000;
   assign mem[9327] = 32'b11111011100110001110100000000000;
   assign mem[9328] = 32'b00000010000110110101000111111100;
   assign mem[9329] = 32'b00000001001100100110001011111100;
   assign mem[9330] = 32'b00000001111100010001010011010010;
   assign mem[9331] = 32'b11110011010100010101110100010000;
   assign mem[9332] = 32'b11111000001010011001111001111000;
   assign mem[9333] = 32'b00000010100110110010001000011000;
   assign mem[9334] = 32'b00000001000001101001010111011000;
   assign mem[9335] = 32'b00000000101101011110111110100111;
   assign mem[9336] = 32'b00000111100000101100110010111000;
   assign mem[9337] = 32'b11111111000111000101101111101000;
   assign mem[9338] = 32'b11111101110110110010100110110000;
   assign mem[9339] = 32'b00000010110100101000110011010100;
   assign mem[9340] = 32'b11111100100100100100000110000000;
   assign mem[9341] = 32'b11111101011110000101001110000000;
   assign mem[9342] = 32'b00000111100011111110000001101000;
   assign mem[9343] = 32'b11110111011100100101110111110000;
   assign mem[9344] = 32'b00001100110110110100110010110000;
   assign mem[9345] = 32'b11111011111110010010111010011000;
   assign mem[9346] = 32'b11110110100010100110101010100000;
   assign mem[9347] = 32'b00000110110101010110110011010000;
   assign mem[9348] = 32'b11111111100001010011111010110000;
   assign mem[9349] = 32'b11111101000011101111010001100000;
   assign mem[9350] = 32'b00000110101110000101100001000000;
   assign mem[9351] = 32'b00000011011010001001000100001000;
   assign mem[9352] = 32'b00000110001010111000111111011000;
   assign mem[9353] = 32'b11111000111011101100011101110000;
   assign mem[9354] = 32'b11101011010000101101010000000000;
   assign mem[9355] = 32'b00001000101000110011011000110000;
   assign mem[9356] = 32'b00000011000110101101000010110000;
   assign mem[9357] = 32'b11101110001111000010111011000000;
   assign mem[9358] = 32'b11111001101100001010110011110000;
   assign mem[9359] = 32'b11110110100010000100100001110000;
   assign mem[9360] = 32'b00000110010101101100100000110000;
   assign mem[9361] = 32'b00000001101100110101111000100010;
   assign mem[9362] = 32'b11111010111010010100010010010000;
   assign mem[9363] = 32'b11111011111111000111101011011000;
   assign mem[9364] = 32'b00000100110100110101000001100000;
   assign mem[9365] = 32'b00000101100001101010010101101000;
   assign mem[9366] = 32'b11111101100100111101011010001000;
   assign mem[9367] = 32'b00001000110000101010011001010000;
   assign mem[9368] = 32'b00000000000011011011100111111011;
   assign mem[9369] = 32'b11111010101100111111000101110000;
   assign mem[9370] = 32'b11110001011011110000101001100000;
   assign mem[9371] = 32'b11111101101011110101100010000100;
   assign mem[9372] = 32'b11110111011110101111101101000000;
   assign mem[9373] = 32'b00000101000001001101000011111000;
   assign mem[9374] = 32'b00000010111011111111000011001000;
   assign mem[9375] = 32'b11111111011111101010100011000100;
   assign mem[9376] = 32'b11111011101010010001111110010000;
   assign mem[9377] = 32'b11111011101111110010111100100000;
   assign mem[9378] = 32'b11111110011101001111011110100000;
   assign mem[9379] = 32'b00000110001001111111110110111000;
   assign mem[9380] = 32'b00000011111001000110011001000100;
   assign mem[9381] = 32'b00001011111100001110000000010000;
   assign mem[9382] = 32'b11110111010100110111010011100000;
   assign mem[9383] = 32'b11111001000111010110110010010000;
   assign mem[9384] = 32'b11111001100110111011101001000000;
   assign mem[9385] = 32'b00001111111010110101100011000000;
   assign mem[9386] = 32'b00000000101000101111011101110011;
   assign mem[9387] = 32'b11110000110110000100010001100000;
   assign mem[9388] = 32'b11111010010000101111001111011000;
   assign mem[9389] = 32'b11111111110110011100101111000001;
   assign mem[9390] = 32'b00000001001010000001100111011110;
   assign mem[9391] = 32'b11111101100011110011001010101000;
   assign mem[9392] = 32'b11111111001100101100011000010010;
   assign mem[9393] = 32'b00000010000101101101001101000100;
   assign mem[9394] = 32'b00000010110001101001100111011000;
   assign mem[9395] = 32'b11111111100011001111101110110011;
   assign mem[9396] = 32'b00000011011011101100001110010000;
   assign mem[9397] = 32'b11111101101111110101010011000000;
   assign mem[9398] = 32'b11111101001100110111110100111000;
   assign mem[9399] = 32'b00000010100111111111101111111000;
   assign mem[9400] = 32'b00001011001000011101001001000000;
   assign mem[9401] = 32'b11111010010111000000110001000000;
   assign mem[9402] = 32'b11111111101110011110000000111001;
   assign mem[9403] = 32'b00000011100111110110000110110100;
   assign mem[9404] = 32'b00000101100010100110110001111000;
   assign mem[9405] = 32'b11111001110101101110110111011000;
   assign mem[9406] = 32'b11111011010101110101111011111000;
   assign mem[9407] = 32'b00000011110101001100010011100000;
   assign mem[9408] = 32'b11111010111001001101001010101000;
   assign mem[9409] = 32'b00000011111010000000111010101100;
   assign mem[9410] = 32'b00000011111111110011100111110000;
   assign mem[9411] = 32'b11110001000001100110110000000000;
   assign mem[9412] = 32'b11111011101010110000010001010000;
   assign mem[9413] = 32'b00000000010001111100111100110100;
   assign mem[9414] = 32'b11110101101110001011011001000000;
   assign mem[9415] = 32'b00000100100101101000111000011000;
   assign mem[9416] = 32'b00000101001101010011000100101000;
   assign mem[9417] = 32'b00000000001011110111011110110011;
   assign mem[9418] = 32'b00000000110100001110011101011000;
   assign mem[9419] = 32'b00000001110001001101011010100010;
   assign mem[9420] = 32'b00001010101101001100100011000000;
   assign mem[9421] = 32'b11111110100010111111011100101110;
   assign mem[9422] = 32'b11110010110110101000111011100000;
   assign mem[9423] = 32'b11111000010111100001111100110000;
   assign mem[9424] = 32'b11110101100111010101110101110000;
   assign mem[9425] = 32'b00001001010110100000101001110000;
   assign mem[9426] = 32'b00000000111011011111101001101100;
   assign mem[9427] = 32'b00001011111011100010011111000000;
   assign mem[9428] = 32'b11111001100000000100101110100000;
   assign mem[9429] = 32'b11100100101100111100010011100000;
   assign mem[9430] = 32'b11111111101110101000110111011000;
   assign mem[9431] = 32'b11111110010110010010101001011000;
   assign mem[9432] = 32'b11111110100011010010000001100000;
   assign mem[9433] = 32'b00000010100101101011001011110100;
   assign mem[9434] = 32'b00000001100000110101000000111000;
   assign mem[9435] = 32'b11111101111111010111000000011100;
   assign mem[9436] = 32'b11111011011111000000010011110000;
   assign mem[9437] = 32'b00000000110111010010110101100010;
   assign mem[9438] = 32'b11111101000000110010111110001100;
   assign mem[9439] = 32'b11111011111110001010110100111000;
   assign mem[9440] = 32'b11111100010010011000100101001000;
   assign mem[9441] = 32'b11111101100101000101100100111000;
   assign mem[9442] = 32'b11111001010001111101100011100000;
   assign mem[9443] = 32'b11111011111100010010100010100000;
   assign mem[9444] = 32'b00000011101011000010011000110000;
   assign mem[9445] = 32'b11110111110010001010100110010000;
   assign mem[9446] = 32'b00000011010011100011101100001100;
   assign mem[9447] = 32'b00001000000011101110000010000000;
   assign mem[9448] = 32'b11111011111100101111110011101000;
   assign mem[9449] = 32'b00000101001110001010111101110000;
   assign mem[9450] = 32'b00000000101100001100010110111010;
   assign mem[9451] = 32'b11111101101000000101001111110000;
   assign mem[9452] = 32'b00001101111101011110111110100000;
   assign mem[9453] = 32'b11110010110101000001110000100000;
   assign mem[9454] = 32'b00000001010100101000111110001010;
   assign mem[9455] = 32'b11110100010010001101010010100000;
   assign mem[9456] = 32'b11111010100111011110101110100000;
   assign mem[9457] = 32'b11110100011101110100111111000000;
   assign mem[9458] = 32'b00001000100110011010010111000000;
   assign mem[9459] = 32'b11111001001010001001000011001000;
   assign mem[9460] = 32'b00000010001000000101011100000000;
   assign mem[9461] = 32'b11110011011000000100000100000000;
   assign mem[9462] = 32'b00000110111011111100110110100000;
   assign mem[9463] = 32'b11111001000111100011110110001000;
   assign mem[9464] = 32'b11111101111010111111001011101100;
   assign mem[9465] = 32'b11101100010011010000100111100000;
   assign mem[9466] = 32'b00000010101100001110011001011100;
   assign mem[9467] = 32'b00000010111010101000101001001100;
   assign mem[9468] = 32'b00001011100111100101101011000000;
   assign mem[9469] = 32'b00000001001011010111111110000100;
   assign mem[9470] = 32'b00010000001011101111111011000000;
   assign mem[9471] = 32'b00000111100011011000010111101000;
   assign mem[9472] = 32'b11111111001010001100011111011100;
   assign mem[9473] = 32'b11101011011010000011101011100000;
   assign mem[9474] = 32'b11110010111100101111010110100000;
   assign mem[9475] = 32'b11111011011011100001111011101000;
   assign mem[9476] = 32'b11111100110001001011011110111100;
   assign mem[9477] = 32'b00000000001100011000000000000011;
   assign mem[9478] = 32'b11111100100110000001000000011000;
   assign mem[9479] = 32'b11111100000011000101001010101100;
   assign mem[9480] = 32'b00000010001011101111000100111000;
   assign mem[9481] = 32'b11110100100011010100000101000000;
   assign mem[9482] = 32'b00000101100010101001111101000000;
   assign mem[9483] = 32'b11111010010111011010000011110000;
   assign mem[9484] = 32'b00000000100101010110101000100100;
   assign mem[9485] = 32'b00000000111000111110111001110110;
   assign mem[9486] = 32'b11111100011111111100000101011100;
   assign mem[9487] = 32'b00000011111100101010101110010100;
   assign mem[9488] = 32'b00000111111100111110110100111000;
   assign mem[9489] = 32'b11110110000111001110001111100000;
   assign mem[9490] = 32'b11110110011100111111110101110000;
   assign mem[9491] = 32'b11110000010011111000011001010000;
   assign mem[9492] = 32'b00000010111010011011101001111100;
   assign mem[9493] = 32'b00000001000100000100111001010100;
   assign mem[9494] = 32'b00000010011000100010011111110000;
   assign mem[9495] = 32'b00000111011111111011100100101000;
   assign mem[9496] = 32'b00000001010100111100000100111100;
   assign mem[9497] = 32'b00000001011101010001001111000000;
   assign mem[9498] = 32'b00000000010101000001101110101101;
   assign mem[9499] = 32'b11110001100110100111111010010000;
   assign mem[9500] = 32'b11111110101100111101101011011100;
   assign mem[9501] = 32'b11111101011011100100110111110000;
   assign mem[9502] = 32'b00000100011010000010001000101000;
   assign mem[9503] = 32'b11111011011000101010011000011000;
   assign mem[9504] = 32'b00000111011011001100000110010000;
   assign mem[9505] = 32'b11111001010110110000110111111000;
   assign mem[9506] = 32'b11110101010010011011100010110000;
   assign mem[9507] = 32'b11111100011110100100100010000000;
   assign mem[9508] = 32'b00001101000111100110010000010000;
   assign mem[9509] = 32'b00000101110000111010000011101000;
   assign mem[9510] = 32'b11111111111000010011001101111111;
   assign mem[9511] = 32'b11110111100101011000111100110000;
   assign mem[9512] = 32'b00000010101011101111010100000000;
   assign mem[9513] = 32'b00000011011110001111100000100100;
   assign mem[9514] = 32'b00000000101110001011010111001010;
   assign mem[9515] = 32'b11111011010100101011101011101000;
   assign mem[9516] = 32'b11110101101000110011110111010000;
   assign mem[9517] = 32'b00000100000001011101001101000000;
   assign mem[9518] = 32'b00000010000111110011101110100000;
   assign mem[9519] = 32'b00000010011000000111110011100000;
   assign mem[9520] = 32'b11111101011111011001001000110000;
   assign mem[9521] = 32'b11111000011100111001011100111000;
   assign mem[9522] = 32'b11111100100111011101100001100000;
   assign mem[9523] = 32'b00000110011010111111001101111000;
   assign mem[9524] = 32'b00000000101110110100011100001101;
   assign mem[9525] = 32'b11111110111110001100101101110010;
   assign mem[9526] = 32'b00000110010001010011011011011000;
   assign mem[9527] = 32'b00000010011001111101101100100000;
   assign mem[9528] = 32'b11111000111011100001010111010000;
   assign mem[9529] = 32'b00000111000001011100111100100000;
   assign mem[9530] = 32'b00000110011111001110010010111000;
   assign mem[9531] = 32'b00000011100001100111101001110000;
   assign mem[9532] = 32'b11110110001000101100001100010000;
   assign mem[9533] = 32'b11111001010011010010010111000000;
   assign mem[9534] = 32'b11110101011011000100101000000000;
   assign mem[9535] = 32'b00001000010111100101111110000000;
   assign mem[9536] = 32'b00000011001010011000111101001000;
   assign mem[9537] = 32'b11111110110000011110011011100010;
   assign mem[9538] = 32'b00000001101011111001110110000110;
   assign mem[9539] = 32'b11111010101110001001010010010000;
   assign mem[9540] = 32'b11111001000001101111100011110000;
   assign mem[9541] = 32'b00000000110010001000110111011110;
   assign mem[9542] = 32'b11111110100110001001011110000110;
   assign mem[9543] = 32'b11111111010110011100101100101110;
   assign mem[9544] = 32'b11111110001110000001010110001110;
   assign mem[9545] = 32'b00000011000100011111000110110100;
   assign mem[9546] = 32'b00000100001100011110000101111000;
   assign mem[9547] = 32'b00000010000110010101001000111000;
   assign mem[9548] = 32'b11110111111111011110101010010000;
   assign mem[9549] = 32'b00000010100111011010111011001100;
   assign mem[9550] = 32'b11111111100010000000101011111011;
   assign mem[9551] = 32'b11111110010101000010011110000110;
   assign mem[9552] = 32'b11111110100010000001001101011010;
   assign mem[9553] = 32'b00000000000010110110001100110101;
   assign mem[9554] = 32'b00000001101010100110001001100000;
   assign mem[9555] = 32'b00000101110000011110110101111000;
   assign mem[9556] = 32'b00000101001111111001011101111000;
   assign mem[9557] = 32'b11111011010100110110110010000000;
   assign mem[9558] = 32'b11110111111010100101101010000000;
   assign mem[9559] = 32'b11111111010010110110001001101110;
   assign mem[9560] = 32'b11111101110010011011110111100100;
   assign mem[9561] = 32'b00000011001001001011110001101100;
   assign mem[9562] = 32'b00001100000001101000110001010000;
   assign mem[9563] = 32'b11110101000010010111110001110000;
   assign mem[9564] = 32'b11111100011010001101011010010000;
   assign mem[9565] = 32'b11111010001000010111111111101000;
   assign mem[9566] = 32'b00000000011111111110001110101010;
   assign mem[9567] = 32'b11110110111111101001111100010000;
   assign mem[9568] = 32'b11111001110011101010000111000000;
   assign mem[9569] = 32'b00000101111111010101100110110000;
   assign mem[9570] = 32'b00000000000110011111100011000100;
   assign mem[9571] = 32'b11111011010001101001000110110000;
   assign mem[9572] = 32'b00000010111000100111110100000100;
   assign mem[9573] = 32'b11110001010000001011110110010000;
   assign mem[9574] = 32'b11111111111111100110010000001110;
   assign mem[9575] = 32'b11110100001110001000101110010000;
   assign mem[9576] = 32'b11111001011101110110110110100000;
   assign mem[9577] = 32'b00000000001101101101100101000100;
   assign mem[9578] = 32'b00000000111010011001110001011110;
   assign mem[9579] = 32'b00000000100011010101111001101000;
   assign mem[9580] = 32'b00001011011110011111011010100000;
   assign mem[9581] = 32'b11111001011111010110100100010000;
   assign mem[9582] = 32'b00001101101111001001101001100000;
   assign mem[9583] = 32'b11100110011000111010110100000000;
   assign mem[9584] = 32'b00001100001011101100011001010000;
   assign mem[9585] = 32'b11110001100100101101111111010000;
   assign mem[9586] = 32'b11110010001100100000101101010000;
   assign mem[9587] = 32'b11111001011101000010000011000000;
   assign mem[9588] = 32'b11110010011011010001110000110000;
   assign mem[9589] = 32'b11111011010001000110101000010000;
   assign mem[9590] = 32'b00000100000110010111110101101000;
   assign mem[9591] = 32'b11110111101100000001101101110000;
   assign mem[9592] = 32'b00001000101010111111111000000000;
   assign mem[9593] = 32'b11101001000011011001111111000000;
   assign mem[9594] = 32'b00000100110000101111000100101000;
   assign mem[9595] = 32'b11110100011010001111001000100000;
   assign mem[9596] = 32'b11111011111011000101011001100000;
   assign mem[9597] = 32'b00000010011101001000000010110100;
   assign mem[9598] = 32'b11111110000001100111101101011010;
   assign mem[9599] = 32'b11111101000000111011111100101100;
   assign mem[9600] = 32'b11111010101101110111000011000000;
   assign mem[9601] = 32'b00001010001000110101000100000000;
   assign mem[9602] = 32'b00000100001001011110101000100000;
   assign mem[9603] = 32'b00000011011001101101110110000100;
   assign mem[9604] = 32'b00000010000010101101101111111000;
   assign mem[9605] = 32'b11111111101101001111001011111000;
   assign mem[9606] = 32'b11111010111110001100100010110000;
   assign mem[9607] = 32'b11111010000110011110110001101000;
   assign mem[9608] = 32'b11111010000000111110011100010000;
   assign mem[9609] = 32'b00000110000110001000011011111000;
   assign mem[9610] = 32'b11111010101001101011111000100000;
   assign mem[9611] = 32'b11111101101011010100101010100100;
   assign mem[9612] = 32'b11111001000101000101010111111000;
   assign mem[9613] = 32'b00001010100100100011011101000000;
   assign mem[9614] = 32'b11111110000110011110101101011010;
   assign mem[9615] = 32'b11111111001111011110101101010010;
   assign mem[9616] = 32'b00000100110001011101111111110000;
   assign mem[9617] = 32'b00000011101010111101010100111000;
   assign mem[9618] = 32'b11111100100100011011110010000000;
   assign mem[9619] = 32'b11111011101001111011001100000000;
   assign mem[9620] = 32'b11111100001111010111100111100000;
   assign mem[9621] = 32'b11101101010110010111011001000000;
   assign mem[9622] = 32'b11110100111110011101000100000000;
   assign mem[9623] = 32'b00000011011000111100011111111000;
   assign mem[9624] = 32'b00000101001000001101001110010000;
   assign mem[9625] = 32'b00000010111110011011111110110000;
   assign mem[9626] = 32'b00000001111011001001001000101100;
   assign mem[9627] = 32'b11110000101111000011110000110000;
   assign mem[9628] = 32'b11111011100100011011111011111000;
   assign mem[9629] = 32'b11111100111111101011010010110100;
   assign mem[9630] = 32'b11111111000011001101010100110001;
   assign mem[9631] = 32'b00000110110000100100101110101000;
   assign mem[9632] = 32'b11110101000011100011111010110000;
   assign mem[9633] = 32'b00000000110110000100101111011001;
   assign mem[9634] = 32'b00001000011101011101111110110000;
   assign mem[9635] = 32'b00000010111011111010100001110100;
   assign mem[9636] = 32'b11110111000001011111101010000000;
   assign mem[9637] = 32'b11111011010100101010101111101000;
   assign mem[9638] = 32'b11110111110000000111110101100000;
   assign mem[9639] = 32'b00000000011010111100001010111011;
   assign mem[9640] = 32'b11110001100101011010001001110000;
   assign mem[9641] = 32'b00000011011010010010111011111000;
   assign mem[9642] = 32'b11111110000000011001001100110110;
   assign mem[9643] = 32'b11111101100101010100111010101000;
   assign mem[9644] = 32'b00000011100100001011011110101100;
   assign mem[9645] = 32'b00000100110000101001011111110000;
   assign mem[9646] = 32'b11101111111001110111000101100000;
   assign mem[9647] = 32'b00000010111101100111010100101000;
   assign mem[9648] = 32'b00000111000011011100000111001000;
   assign mem[9649] = 32'b11111010010101101111111000110000;
   assign mem[9650] = 32'b00000100011000101100000001101000;
   assign mem[9651] = 32'b11101101101010001001001010000000;
   assign mem[9652] = 32'b00000110101101100001110011011000;
   assign mem[9653] = 32'b11111000101110111011111111101000;
   assign mem[9654] = 32'b11111111010011110000001111101011;
   assign mem[9655] = 32'b00000000001110100101110101110111;
   assign mem[9656] = 32'b11111011101010111100111111111000;
   assign mem[9657] = 32'b11111101111111010000110010101100;
   assign mem[9658] = 32'b00000001000101011101101100001110;
   assign mem[9659] = 32'b00000010010110100111001100011100;
   assign mem[9660] = 32'b00000100110000011011101011111000;
   assign mem[9661] = 32'b00000001101100101111001101001110;
   assign mem[9662] = 32'b00000110010000001101000100101000;
   assign mem[9663] = 32'b11111011111000011101001110100000;
   assign mem[9664] = 32'b11110111110011110110011111110000;
   assign mem[9665] = 32'b11110011100010111001000011010000;
   assign mem[9666] = 32'b11111111110111010100010101001101;
   assign mem[9667] = 32'b00001000001100111001101010010000;
   assign mem[9668] = 32'b11111011001000001100000101011000;
   assign mem[9669] = 32'b00000101000101111000111010100000;
   assign mem[9670] = 32'b00000001111011100101110011100010;
   assign mem[9671] = 32'b00001001001001011100010010100000;
   assign mem[9672] = 32'b11111011101111001010010001000000;
   assign mem[9673] = 32'b11110111110011110010101001110000;
   assign mem[9674] = 32'b00000010101110011011100101100100;
   assign mem[9675] = 32'b00000011111101111110100010000100;
   assign mem[9676] = 32'b11111101111111010011011100110100;
   assign mem[9677] = 32'b00000110111110010100110111001000;
   assign mem[9678] = 32'b11111111000100000011011110011101;
   assign mem[9679] = 32'b11110111110100101011000110100000;
   assign mem[9680] = 32'b11101010100101100010111000100000;
   assign mem[9681] = 32'b00000111000001110101010010111000;
   assign mem[9682] = 32'b11111111001011001101010010100100;
   assign mem[9683] = 32'b00000111001100100010000001001000;
   assign mem[9684] = 32'b11111111001011011001000010101110;
   assign mem[9685] = 32'b00001000010101000100111010010000;
   assign mem[9686] = 32'b11101110011110001000110000100000;
   assign mem[9687] = 32'b11111011111010100000011100011000;
   assign mem[9688] = 32'b00000011011111101110001101101000;
   assign mem[9689] = 32'b11111111001111011100110000011011;
   assign mem[9690] = 32'b00000100110110100111111111010000;
   assign mem[9691] = 32'b11111101000001010011111110001100;
   assign mem[9692] = 32'b00000001101010110000010101110100;
   assign mem[9693] = 32'b11111001010101110101111111000000;
   assign mem[9694] = 32'b11111110000011111000110001010000;
   assign mem[9695] = 32'b00000010011011010000001010000000;
   assign mem[9696] = 32'b00000010010110110001010010001000;
   assign mem[9697] = 32'b11110111101111010001001001010000;
   assign mem[9698] = 32'b00000010000000111011010000101000;
   assign mem[9699] = 32'b11111111000110111110011001011010;
   assign mem[9700] = 32'b11111100110000111001010110101100;
   assign mem[9701] = 32'b00000000011110001101000000010010;
   assign mem[9702] = 32'b00000011110100000110100111110100;
   assign mem[9703] = 32'b11111101011000100110101110110100;
   assign mem[9704] = 32'b00000001000011110010111010101110;
   assign mem[9705] = 32'b00000110010011110100111001010000;
   assign mem[9706] = 32'b11111011111100100111001100101000;
   assign mem[9707] = 32'b00000000100100000010101100110011;
   assign mem[9708] = 32'b11111011101111001111000001000000;
   assign mem[9709] = 32'b11110000111000010010001101010000;
   assign mem[9710] = 32'b00000101111001110000011001101000;
   assign mem[9711] = 32'b11111011000000110110000011101000;
   assign mem[9712] = 32'b11111011011101101101010011010000;
   assign mem[9713] = 32'b11111101101110110101000010001100;
   assign mem[9714] = 32'b00000001000101111101101110010100;
   assign mem[9715] = 32'b11111111110000110100001111000100;
   assign mem[9716] = 32'b00000110001011000010111011110000;
   assign mem[9717] = 32'b11111011101010011110001100111000;
   assign mem[9718] = 32'b00000011111110101101111011110100;
   assign mem[9719] = 32'b11111111111110010111100100110100;
   assign mem[9720] = 32'b11111010100000101100100011110000;
   assign mem[9721] = 32'b00000111010111110001101000010000;
   assign mem[9722] = 32'b11111111111000110110000010010010;
   assign mem[9723] = 32'b00000010100001011111010010110100;
   assign mem[9724] = 32'b11111011010100111010010011110000;
   assign mem[9725] = 32'b11111110110101101010101011110110;
   assign mem[9726] = 32'b11111110011101100010111000010000;
   assign mem[9727] = 32'b11111111001011100010010100100100;
   assign mem[9728] = 32'b11111000110101001000011101000000;
   assign mem[9729] = 32'b00000001000001100000110000010000;
   assign mem[9730] = 32'b11111011010010001101010100001000;
   assign mem[9731] = 32'b00000100000011010111101101100000;
   assign mem[9732] = 32'b11111110011001001100000100010010;
   assign mem[9733] = 32'b00000111000011001000001000000000;
   assign mem[9734] = 32'b11101110101101010010011010100000;
   assign mem[9735] = 32'b00000011011000001001110111100000;
   assign mem[9736] = 32'b11110011110001100101100110000000;
   assign mem[9737] = 32'b11110111111101010011011100010000;
   assign mem[9738] = 32'b11111011001010001010000011100000;
   assign mem[9739] = 32'b00000010001111001101010000100000;
   assign mem[9740] = 32'b00000111000111100111011110000000;
   assign mem[9741] = 32'b11111111011101001010111100000110;
   assign mem[9742] = 32'b00000011111101000000011110101100;
   assign mem[9743] = 32'b11111111000001100110011011001111;
   assign mem[9744] = 32'b00000111001101100001111100001000;
   assign mem[9745] = 32'b11111100100100001100100111110000;
   assign mem[9746] = 32'b11111110111110100000101011111110;
   assign mem[9747] = 32'b11110011000100011111110100110000;
   assign mem[9748] = 32'b11110110100000111101010001010000;
   assign mem[9749] = 32'b11111100000110010110111100011100;
   assign mem[9750] = 32'b00000110000101011110001001111000;
   assign mem[9751] = 32'b11111001100100000011101111110000;
   assign mem[9752] = 32'b00000000011011110011100010100000;
   assign mem[9753] = 32'b11111010110010000010110110010000;
   assign mem[9754] = 32'b11111110001011011011001101011100;
   assign mem[9755] = 32'b11111010100111100010001010110000;
   assign mem[9756] = 32'b00000011001010010001000000010100;
   assign mem[9757] = 32'b11111101011111100111000001100100;
   assign mem[9758] = 32'b00000110111111110110100110011000;
   assign mem[9759] = 32'b11111011000010110101001010111000;
   assign mem[9760] = 32'b11111011101000001100110101101000;
   assign mem[9761] = 32'b00001000001010000101111000100000;
   assign mem[9762] = 32'b00000010011000100000010011001100;
   assign mem[9763] = 32'b11111110001110001010001000001000;
   assign mem[9764] = 32'b00000110101010101100111000000000;
   assign mem[9765] = 32'b00000000111110001101010110111011;
   assign mem[9766] = 32'b11111100110111000011101001100100;
   assign mem[9767] = 32'b11111110111011100001000001010110;
   assign mem[9768] = 32'b11111000100001010111110011011000;
   assign mem[9769] = 32'b11111010100100000110100000100000;
   assign mem[9770] = 32'b00000000011000000100000111110010;
   assign mem[9771] = 32'b11110110010001100011100010010000;
   assign mem[9772] = 32'b00000000100100101100100101010010;
   assign mem[9773] = 32'b00000010001101110101110011001100;
   assign mem[9774] = 32'b00000001110110011011111001111100;
   assign mem[9775] = 32'b11111011101110101100110000101000;
   assign mem[9776] = 32'b00000100100101111100110101011000;
   assign mem[9777] = 32'b11111101010111100111001111101100;
   assign mem[9778] = 32'b11111100110101111101111001010000;
   assign mem[9779] = 32'b11111011101011100000000000001000;
   assign mem[9780] = 32'b11111001010001001100010110100000;
   assign mem[9781] = 32'b11110111110010010011101011000000;
   assign mem[9782] = 32'b11110110110110110101000000000000;
   assign mem[9783] = 32'b00000001011101011101101100001010;
   assign mem[9784] = 32'b00001111001001111010100111000000;
   assign mem[9785] = 32'b00000011011110110100101100111100;
   assign mem[9786] = 32'b11110000111111011011111011100000;
   assign mem[9787] = 32'b00000101100011100011110010101000;
   assign mem[9788] = 32'b00000100100010001110000100001000;
   assign mem[9789] = 32'b11111110001110110101111011000100;
   assign mem[9790] = 32'b11111110101000110000110100000110;
   assign mem[9791] = 32'b00000110100010111101111001101000;
   assign mem[9792] = 32'b00001100000000000011010010100000;
   assign mem[9793] = 32'b11111101100010111110010001111000;
   assign mem[9794] = 32'b11110101011100001110100111100000;
   assign mem[9795] = 32'b11111101010101001110100011111100;
   assign mem[9796] = 32'b11111110010011000100011111101000;
   assign mem[9797] = 32'b00001011100110011011010101110000;
   assign mem[9798] = 32'b00000001000110100010000010111110;
   assign mem[9799] = 32'b11100111000000010111010010100000;
   assign mem[9800] = 32'b00000011011100101110110101111000;
   assign mem[9801] = 32'b11110110011000011001110000110000;
   assign mem[9802] = 32'b00000001010101110111110000001110;
   assign mem[9803] = 32'b11111001011101110000111001101000;
   assign mem[9804] = 32'b00000011111110000110011110010100;
   assign mem[9805] = 32'b11110011101100110101111010110000;
   assign mem[9806] = 32'b00000100010101100001100001001000;
   assign mem[9807] = 32'b00000100010110000111000101111000;
   assign mem[9808] = 32'b11111110011010001001100000001010;
   assign mem[9809] = 32'b00000111111101100011010111101000;
   assign mem[9810] = 32'b11110010011010101110111010010000;
   assign mem[9811] = 32'b00000010110001010000110001101000;
   assign mem[9812] = 32'b00000101101011100110111100000000;
   assign mem[9813] = 32'b11111000111011101110101101010000;
   assign mem[9814] = 32'b11111100011010001001100100000000;
   assign mem[9815] = 32'b11111011001000010111011101010000;
   assign mem[9816] = 32'b11111001100111010001100111000000;
   assign mem[9817] = 32'b00000001010011100010110101111110;
   assign mem[9818] = 32'b00000100000010010101000110000000;
   assign mem[9819] = 32'b11111010001001111001100101000000;
   assign mem[9820] = 32'b00001010011101010110010110010000;
   assign mem[9821] = 32'b11111101010110101110101100101000;
   assign mem[9822] = 32'b11111111111100011010000011010011;
   assign mem[9823] = 32'b11110010101010111000010011100000;
   assign mem[9824] = 32'b00000101011111000111000101101000;
   assign mem[9825] = 32'b11111111110010010000100011000111;
   assign mem[9826] = 32'b00000000100111101010001001011111;
   assign mem[9827] = 32'b00000111111001011000111000111000;
   assign mem[9828] = 32'b11111111101000110110011010111111;
   assign mem[9829] = 32'b11111001100000000010100101110000;
   assign mem[9830] = 32'b00000010110000101100111010010000;
   assign mem[9831] = 32'b11110011000000111010001011110000;
   assign mem[9832] = 32'b11111110111001000000111010000000;
   assign mem[9833] = 32'b00000101000111100000011011111000;
   assign mem[9834] = 32'b00000001010001010111001111001100;
   assign mem[9835] = 32'b11111111000111000100110010110110;
   assign mem[9836] = 32'b00000110001111111111101100011000;
   assign mem[9837] = 32'b11111010101010011111100001111000;
   assign mem[9838] = 32'b11111100110000011101110110010100;
   assign mem[9839] = 32'b11111101101011011110100100001000;
   assign mem[9840] = 32'b00000100101000001011001001111000;
   assign mem[9841] = 32'b11110000111001111011001010010000;
   assign mem[9842] = 32'b11111010111100011110000111000000;
   assign mem[9843] = 32'b00000101101010001011010100011000;
   assign mem[9844] = 32'b11111101011111100101000010000000;
   assign mem[9845] = 32'b00000011100001100111101011000100;
   assign mem[9846] = 32'b00000101100000010101111001000000;
   assign mem[9847] = 32'b11111011100011010111000100010000;
   assign mem[9848] = 32'b11111101000100011010011001010000;
   assign mem[9849] = 32'b00000000011000100110000001110010;
   assign mem[9850] = 32'b00000001111000100010011001111000;
   assign mem[9851] = 32'b00001011010010011011001110010000;
   assign mem[9852] = 32'b11111000111011010100101101010000;
   assign mem[9853] = 32'b00000011000100100000011010111000;
   assign mem[9854] = 32'b11111101110001010010000101111000;
   assign mem[9855] = 32'b11110001101110011110100010000000;
   assign mem[9856] = 32'b11111001101010000111111001011000;
   assign mem[9857] = 32'b00001011011000111111111011000000;
   assign mem[9858] = 32'b11110110011010010011001010110000;
   assign mem[9859] = 32'b11111100000011110010100001110100;
   assign mem[9860] = 32'b00000101110111100100001110010000;
   assign mem[9861] = 32'b11101011111001101000110011100000;
   assign mem[9862] = 32'b11110110111110111101000000110000;
   assign mem[9863] = 32'b00000000100000101010110000101110;
   assign mem[9864] = 32'b11111000111110101011111111000000;
   assign mem[9865] = 32'b11110000101000111001000110000000;
   assign mem[9866] = 32'b00000001011001110110110011101010;
   assign mem[9867] = 32'b11111110000101011001111110110000;
   assign mem[9868] = 32'b11111011011101000010101001110000;
   assign mem[9869] = 32'b00001000101010100000010111100000;
   assign mem[9870] = 32'b11111011101101011110011001001000;
   assign mem[9871] = 32'b00000001010100000010110001101110;
   assign mem[9872] = 32'b00000100100100110101000111110000;
   assign mem[9873] = 32'b11111001101010001001000111010000;
   assign mem[9874] = 32'b11111101000011101110110101001000;
   assign mem[9875] = 32'b11111111001011110100101010011001;
   assign mem[9876] = 32'b11111101101110011010010000010000;
   assign mem[9877] = 32'b11111110100001111110010010110010;
   assign mem[9878] = 32'b00000101111100000111101000100000;
   assign mem[9879] = 32'b11110111000101100011100110100000;
   assign mem[9880] = 32'b11111100010100100111101101010100;
   assign mem[9881] = 32'b11111111101011000100010100000001;
   assign mem[9882] = 32'b00001100111100010101110111100000;
   assign mem[9883] = 32'b11111100000110000000110011111100;
   assign mem[9884] = 32'b00000001111001001011100001101100;
   assign mem[9885] = 32'b11111101100001000010000110011000;
   assign mem[9886] = 32'b11111110000101001101011001111010;
   assign mem[9887] = 32'b11110100111100001000110000010000;
   assign mem[9888] = 32'b11111010001001001111000100011000;
   assign mem[9889] = 32'b11111111011010010001010100100010;
   assign mem[9890] = 32'b11101101000001011000101010000000;
   assign mem[9891] = 32'b00000110101100101111011001011000;
   assign mem[9892] = 32'b00000100111110011111000100111000;
   assign mem[9893] = 32'b00000011101011110011101100010100;
   assign mem[9894] = 32'b11110100100010000110010100100000;
   assign mem[9895] = 32'b00000111011111000010101000111000;
   assign mem[9896] = 32'b11110101100100001100100001000000;
   assign mem[9897] = 32'b11111111011111001101100000010010;
   assign mem[9898] = 32'b11111100101010100001101101110100;
   assign mem[9899] = 32'b11111010110110111111100000001000;
   assign mem[9900] = 32'b00000001011110101110000010100000;
   assign mem[9901] = 32'b11101101111110110010010100100000;
   assign mem[9902] = 32'b11111101110101100010000000010100;
   assign mem[9903] = 32'b11111101001111101100110111001100;
   assign mem[9904] = 32'b11111101001100110111010000011000;
   assign mem[9905] = 32'b11111101111111010100000111011100;
   assign mem[9906] = 32'b00000101010110000111000101011000;
   assign mem[9907] = 32'b00001001011001010011001010000000;
   assign mem[9908] = 32'b11111100100010001111000001111100;
   assign mem[9909] = 32'b00000010000111001110100011000000;
   assign mem[9910] = 32'b11111111011011000000001111100111;
   assign mem[9911] = 32'b00000100100010110111101001111000;
   assign mem[9912] = 32'b11111101010101011000100000000000;
   assign mem[9913] = 32'b11111011010000101010001100110000;
   assign mem[9914] = 32'b00000001011101010101110011111100;
   assign mem[9915] = 32'b00000100111101001101110000001000;
   assign mem[9916] = 32'b00000001001010110001000001010010;
   assign mem[9917] = 32'b11111011010111110101110010000000;
   assign mem[9918] = 32'b00000000111011010101001110010100;
   assign mem[9919] = 32'b11111110110100110101011111111000;
   assign mem[9920] = 32'b00001000001100100001010010110000;
   assign mem[9921] = 32'b11110101101000001110011011100000;
   assign mem[9922] = 32'b00000111011110000111111001100000;
   assign mem[9923] = 32'b11110011000011000101000001110000;
   assign mem[9924] = 32'b00000011110110011011011001111000;
   assign mem[9925] = 32'b00000000000011011001001110000011;
   assign mem[9926] = 32'b00000001101001110110111010110000;
   assign mem[9927] = 32'b11110111111000001110010110110000;
   assign mem[9928] = 32'b00000111110111010011010101001000;
   assign mem[9929] = 32'b11110011000111110100111001010000;
   assign mem[9930] = 32'b00000100111010111111111000101000;
   assign mem[9931] = 32'b11101011010100000010100110100000;
   assign mem[9932] = 32'b11111111100011000111010100101001;
   assign mem[9933] = 32'b11110000100010010110001001100000;
   assign mem[9934] = 32'b00000100010100111100111010100000;
   assign mem[9935] = 32'b11111111000011011100001101001101;
   assign mem[9936] = 32'b00000000011100111000111011001100;
   assign mem[9937] = 32'b11111000011101010111101011100000;
   assign mem[9938] = 32'b00000000011110010101101110111100;
   assign mem[9939] = 32'b00001000000100000110101011010000;
   assign mem[9940] = 32'b00000100101101010010100010010000;
   assign mem[9941] = 32'b00000110100010010100001011100000;
   assign mem[9942] = 32'b11111101110010110011001011111000;
   assign mem[9943] = 32'b11111011111100000000010001010000;
   assign mem[9944] = 32'b00000111001010111101101010011000;
   assign mem[9945] = 32'b11110111110101000110110101000000;
   assign mem[9946] = 32'b00000001011100000110111011110010;
   assign mem[9947] = 32'b00000001100100101001001001001010;
   assign mem[9948] = 32'b00000110110010000111100110100000;
   assign mem[9949] = 32'b00000000110000011000000000011111;
   assign mem[9950] = 32'b11110001010010011001011110100000;
   assign mem[9951] = 32'b00000110100110000101110010000000;
   assign mem[9952] = 32'b00000110100111000000000000010000;
   assign mem[9953] = 32'b11111100001001110100000001001000;
   assign mem[9954] = 32'b11111011110011001101111000001000;
   assign mem[9955] = 32'b00000000111110110101010111100111;
   assign mem[9956] = 32'b11111000110100011101100000100000;
   assign mem[9957] = 32'b00000001110011000110101010001000;
   assign mem[9958] = 32'b00001000010100110000101111100000;
   assign mem[9959] = 32'b11110110111101111000001110000000;
   assign mem[9960] = 32'b11111001010011010101011010100000;
   assign mem[9961] = 32'b00000101111111110110111011011000;
   assign mem[9962] = 32'b11110110001100101001100000010000;
   assign mem[9963] = 32'b00000010110100011010001110000000;
   assign mem[9964] = 32'b00000010011011110111110011010100;
   assign mem[9965] = 32'b00000110011010110011110111111000;
   assign mem[9966] = 32'b11101000001111001010100100100000;
   assign mem[9967] = 32'b11111101111110100110010100011000;
   assign mem[9968] = 32'b00000001011100001001011100101100;
   assign mem[9969] = 32'b11111010011111100111011010111000;
   assign mem[9970] = 32'b11111011010101001101111101101000;
   assign mem[9971] = 32'b11111000111101000010001100110000;
   assign mem[9972] = 32'b00000010010111111110000001101000;
   assign mem[9973] = 32'b00000111000001010001011100011000;
   assign mem[9974] = 32'b11110011100011101110100011010000;
   assign mem[9975] = 32'b00001010000001100011010010100000;
   assign mem[9976] = 32'b11110010001100001010101001110000;
   assign mem[9977] = 32'b11110101000001110110011110010000;
   assign mem[9978] = 32'b11111010110001000110001001101000;
   assign mem[9979] = 32'b11111011001101011001000011001000;
   assign mem[9980] = 32'b11111101011101010111101001000100;
   assign mem[9981] = 32'b11111100110110000110001110010100;
   assign mem[9982] = 32'b00000110110101011010101000000000;
   assign mem[9983] = 32'b00000000101100101111001111011100;
   assign mem[9984] = 32'b00000101110000111010101000100000;
   assign mem[9985] = 32'b11111001111011101001110110010000;
   assign mem[9986] = 32'b00000000111001100011000010100110;
   assign mem[9987] = 32'b11110100111011001101010111110000;
   assign mem[9988] = 32'b11111001101101010110100100010000;
   assign mem[9989] = 32'b00000010010110111110011111101100;
   assign mem[9990] = 32'b11101110011000011001010001100000;
   assign mem[9991] = 32'b00000111010011110001110110101000;
   assign mem[9992] = 32'b11111111101100010101101010010100;
   assign mem[9993] = 32'b00000001001101000001111011101000;
   assign mem[9994] = 32'b00000001001100101111001101111010;
   assign mem[9995] = 32'b00000010011100111010101000101000;
   assign mem[9996] = 32'b11101100010101110010010110000000;
   assign mem[9997] = 32'b00000101100011011111001111101000;
   assign mem[9998] = 32'b11111111000000110111000001001001;
   assign mem[9999] = 32'b11111011111010101010110000010000;
   assign mem[10000] = 32'b00000011010011011101010010010100;
   assign mem[10001] = 32'b11101101101000000010100010100000;
   assign mem[10002] = 32'b11111011110010100101100001000000;
   assign mem[10003] = 32'b11110111101110010110001000110000;
   assign mem[10004] = 32'b00000101101110000101100100101000;
   assign mem[10005] = 32'b11111011101101010011010110000000;
   assign mem[10006] = 32'b00000100110010000110100101010000;
   assign mem[10007] = 32'b11111000100110110011110110000000;
   assign mem[10008] = 32'b00000011100011111000000001101000;
   assign mem[10009] = 32'b00000100101100010011011011100000;
   assign mem[10010] = 32'b11111101010110010101100011010000;
   assign mem[10011] = 32'b00000100010101010111110000011000;
   assign mem[10012] = 32'b11111001101101100111011010111000;
   assign mem[10013] = 32'b11111110100100100110001110010100;
   assign mem[10014] = 32'b00000010101111010110011101011100;
   assign mem[10015] = 32'b00000101010011010000001110100000;
   assign mem[10016] = 32'b11110011100111000010011000110000;
   assign mem[10017] = 32'b00000100101001100110110110110000;
   assign mem[10018] = 32'b11111011011100001011001101011000;
   assign mem[10019] = 32'b11111011101001111111100100110000;
   assign mem[10020] = 32'b11111100010111010001110010000100;
   assign mem[10021] = 32'b00000000010100011001110101000010;
   assign mem[10022] = 32'b11111100000000000000011110010100;
   assign mem[10023] = 32'b11111101000111101110100101011100;
   assign mem[10024] = 32'b00000010110001111011000010100100;
   assign mem[10025] = 32'b11111101101101110111100101110100;
   assign mem[10026] = 32'b11111110101000010110101010110000;
   assign mem[10027] = 32'b11111110000011010100110000000000;
   assign mem[10028] = 32'b00000000010111001110000000000111;
   assign mem[10029] = 32'b00000010011110101001010010001100;
   assign mem[10030] = 32'b11111011111111000001111101110000;
   assign mem[10031] = 32'b11111110101111110001001011100100;
   assign mem[10032] = 32'b00000010111001101000111101111100;
   assign mem[10033] = 32'b00000111101010000100010111100000;
   assign mem[10034] = 32'b00000100011001111110001100101000;
   assign mem[10035] = 32'b11111000000111101101111000101000;
   assign mem[10036] = 32'b11111011111111011111111110110000;
   assign mem[10037] = 32'b11110101101011111000000001010000;
   assign mem[10038] = 32'b11111110101110011110011100100100;
   assign mem[10039] = 32'b00000100010111101010000111001000;
   assign mem[10040] = 32'b00000100011111001101111110100000;
   assign mem[10041] = 32'b11111000100001111011101000100000;
   assign mem[10042] = 32'b00000110111111110010010100110000;
   assign mem[10043] = 32'b11111100110100101011001111010100;
   assign mem[10044] = 32'b11111110001010101010100101101000;
   assign mem[10045] = 32'b11110011111001011000101101010000;
   assign mem[10046] = 32'b00000100001110001101111100111000;
   assign mem[10047] = 32'b11110101001110001010100010100000;
   assign mem[10048] = 32'b00000111001011000100100101011000;
   assign mem[10049] = 32'b00000001101101100000010001010110;
   assign mem[10050] = 32'b00000011001100001001110110010100;
   assign mem[10051] = 32'b11111101110011110111000010001100;
   assign mem[10052] = 32'b00000100001101110110110111010000;
   assign mem[10053] = 32'b00000011001010101101010011010000;
   assign mem[10054] = 32'b11111100001111100110100010000000;
   assign mem[10055] = 32'b00000010110001110000110110110000;
   assign mem[10056] = 32'b11111011000010100101100110101000;
   assign mem[10057] = 32'b11111011100100001110001110010000;
   assign mem[10058] = 32'b00000101100111111010010000111000;
   assign mem[10059] = 32'b11111011101000000110111000111000;
   assign mem[10060] = 32'b00000100110001010011101001101000;
   assign mem[10061] = 32'b11111000000000010010001101000000;
   assign mem[10062] = 32'b00000010010011001001101100010100;
   assign mem[10063] = 32'b11110111110110100000000000110000;
   assign mem[10064] = 32'b11111100100110000101010011101100;
   assign mem[10065] = 32'b11111011111110011000101110101000;
   assign mem[10066] = 32'b00001001000110100101011001110000;
   assign mem[10067] = 32'b11110010110101101100101101010000;
   assign mem[10068] = 32'b00000000010010000101110001001011;
   assign mem[10069] = 32'b00000011111100111110011100110100;
   assign mem[10070] = 32'b11111111000101000101110001011010;
   assign mem[10071] = 32'b11111101111101010100000010111000;
   assign mem[10072] = 32'b00000000000111000001010000011000;
   assign mem[10073] = 32'b11111100111001011001101001100100;
   assign mem[10074] = 32'b11111100000111001110111100111100;
   assign mem[10075] = 32'b11111101110100000001000100100000;
   assign mem[10076] = 32'b00000001011010101010111000010010;
   assign mem[10077] = 32'b00000001000111000100011011100110;
   assign mem[10078] = 32'b00000011000101001001001010001100;
   assign mem[10079] = 32'b00000010010101000000001101110100;
   assign mem[10080] = 32'b00000001101011000101001011000010;
   assign mem[10081] = 32'b11110111110101000001110101000000;
   assign mem[10082] = 32'b11111110000011111101011101010010;
   assign mem[10083] = 32'b11111101010110110100011111100000;
   assign mem[10084] = 32'b00000011100100101010110000001000;
   assign mem[10085] = 32'b11111100110111100101000111110100;
   assign mem[10086] = 32'b00000000011101010101111100000000;
   assign mem[10087] = 32'b11111101010001100000110110010000;
   assign mem[10088] = 32'b11111110101111110000011011101100;
   assign mem[10089] = 32'b11111101111111000111001111001000;
   assign mem[10090] = 32'b00000011110111111011010100101100;
   assign mem[10091] = 32'b11111011110111000100111110011000;
   assign mem[10092] = 32'b00000010101101100101111111011000;
   assign mem[10093] = 32'b11110110111010010110100000010000;
   assign mem[10094] = 32'b00000001111000000001110011000100;
   assign mem[10095] = 32'b11111010111111110010010111000000;
   assign mem[10096] = 32'b00000100011010001110010110100000;
   assign mem[10097] = 32'b11111010111111101110010000101000;
   assign mem[10098] = 32'b00000010000010000100100111101000;
   assign mem[10099] = 32'b11110110110101110011010010100000;
   assign mem[10100] = 32'b00001001111111111001010001010000;
   assign mem[10101] = 32'b11111110011011110000001111010000;
   assign mem[10102] = 32'b00000001101010111111010100000100;
   assign mem[10103] = 32'b11101111011010011101001101100000;
   assign mem[10104] = 32'b00000111111010100100111000101000;
   assign mem[10105] = 32'b00000001101100101101100000110110;
   assign mem[10106] = 32'b11111111101000111000010000110101;
   assign mem[10107] = 32'b11111011010110001110100011001000;
   assign mem[10108] = 32'b00000110110010110101100011100000;
   assign mem[10109] = 32'b11111011001101110010000001111000;
   assign mem[10110] = 32'b00000001010100110111010011010110;
   assign mem[10111] = 32'b11111110010100111100001101000010;
   assign mem[10112] = 32'b11111101010010111101110100010100;
   assign mem[10113] = 32'b11111111101111100110000010100100;
   assign mem[10114] = 32'b11111101100110101110010000111000;
   assign mem[10115] = 32'b00000001010100001011101001110100;
   assign mem[10116] = 32'b00000001101000001100111111000000;
   assign mem[10117] = 32'b00000010011110111000001101110000;
   assign mem[10118] = 32'b00000010110101001010000010011100;
   assign mem[10119] = 32'b00000010000111100001110111110100;
   assign mem[10120] = 32'b00000100010111001010110101101000;
   assign mem[10121] = 32'b00000111000111110001101000011000;
   assign mem[10122] = 32'b11111110001100001001100011001000;
   assign mem[10123] = 32'b11111001001001111111111011001000;
   assign mem[10124] = 32'b00000101101001001000110011100000;
   assign mem[10125] = 32'b11111100100010001111010000000100;
   assign mem[10126] = 32'b11111000101011101000100101110000;
   assign mem[10127] = 32'b11111100111001011110010111011000;
   assign mem[10128] = 32'b11111101011111101111111010101100;
   assign mem[10129] = 32'b00000001100101001111100010110100;
   assign mem[10130] = 32'b00000010011011010010010010100000;
   assign mem[10131] = 32'b00000011111011000000001110100100;
   assign mem[10132] = 32'b11111101011100000001011011000100;
   assign mem[10133] = 32'b11111111000001000111010001110111;
   assign mem[10134] = 32'b11111110101111011101011101000010;
   assign mem[10135] = 32'b11111111110101110110001011001101;
   assign mem[10136] = 32'b11111010011011010001101011111000;
   assign mem[10137] = 32'b11111010000011000110100011001000;
   assign mem[10138] = 32'b11111011100010101000110011100000;
   assign mem[10139] = 32'b00000100100101000001000111011000;
   assign mem[10140] = 32'b00000010010010101001000000100100;
   assign mem[10141] = 32'b11111001110110110100011011001000;
   assign mem[10142] = 32'b00000100101100000010110010110000;
   assign mem[10143] = 32'b11110111100110010000000000100000;
   assign mem[10144] = 32'b00000100111100000111100000110000;
   assign mem[10145] = 32'b00000011111010011001010110011000;
   assign mem[10146] = 32'b11111100010011001010101011011100;
   assign mem[10147] = 32'b00000000010111111001011110001101;
   assign mem[10148] = 32'b00000001101010010001010101110010;
   assign mem[10149] = 32'b11111110100011001010001101001110;
   assign mem[10150] = 32'b11111110100000100001010101101110;
   assign mem[10151] = 32'b11111010101100110100011100001000;
   assign mem[10152] = 32'b00001001100001011101010101110000;
   assign mem[10153] = 32'b11111111001100111100101110001000;
   assign mem[10154] = 32'b00000001100001100111100001010100;
   assign mem[10155] = 32'b11111110001101010110011010101010;
   assign mem[10156] = 32'b11111110010000011100000001010100;
   assign mem[10157] = 32'b11111100110111010010101110100100;
   assign mem[10158] = 32'b00000011101011011101011111101000;
   assign mem[10159] = 32'b00000000000101110000010010010111;
   assign mem[10160] = 32'b00000010101010001011001000010100;
   assign mem[10161] = 32'b11111110110010001100010101001000;
   assign mem[10162] = 32'b00000110101101001111110010111000;
   assign mem[10163] = 32'b11111110100011110001011111111100;
   assign mem[10164] = 32'b11111111001100011000111010110111;
   assign mem[10165] = 32'b11111011011010000011111011100000;
   assign mem[10166] = 32'b11111110011000010110000100010110;
   assign mem[10167] = 32'b11111010110111100111001111111000;
   assign mem[10168] = 32'b00000000111010001111110010111111;
   assign mem[10169] = 32'b11111110010001111001110110111000;
   assign mem[10170] = 32'b00000100011000001000010011101000;
   assign mem[10171] = 32'b11111011101001110011011001000000;
   assign mem[10172] = 32'b11111000101100101010011100011000;
   assign mem[10173] = 32'b11111010101100001111111001111000;
   assign mem[10174] = 32'b00000111010111101000011001100000;
   assign mem[10175] = 32'b11111101011101001001101100001000;
   assign mem[10176] = 32'b00000101111111101101010100110000;
   assign mem[10177] = 32'b11110100101100011001110100110000;
   assign mem[10178] = 32'b00000011011100000111001011111000;
   assign mem[10179] = 32'b00000110001001111110111100010000;
   assign mem[10180] = 32'b11111000011011110001000111101000;
   assign mem[10181] = 32'b00000110100100111001110110100000;
   assign mem[10182] = 32'b11111100011000011111000001000000;
   assign mem[10183] = 32'b00000111101011111100011111100000;
   assign mem[10184] = 32'b11111010110010011010110010101000;
   assign mem[10185] = 32'b00000101001011000110011111110000;
   assign mem[10186] = 32'b11110001011010111101101011110000;
   assign mem[10187] = 32'b11110111010111011111101100110000;
   assign mem[10188] = 32'b00000000001001110100100010101110;
   assign mem[10189] = 32'b11110100101110110010110111010000;
   assign mem[10190] = 32'b00000000100101010000001011101011;
   assign mem[10191] = 32'b11111011100100010011110101101000;
   assign mem[10192] = 32'b00000100101011110101110110011000;
   assign mem[10193] = 32'b00000110101011100011111100000000;
   assign mem[10194] = 32'b11110110100110110110010100010000;
   assign mem[10195] = 32'b00000001101011110010101000010100;
   assign mem[10196] = 32'b11110110101011101001110111000000;
   assign mem[10197] = 32'b11111010000100110001110011100000;
   assign mem[10198] = 32'b00000101111001100110001000010000;
   assign mem[10199] = 32'b11101100111010101100101100100000;
   assign mem[10200] = 32'b11101111100101100001011111100000;
   assign mem[10201] = 32'b00000100101110110100001001000000;
   assign mem[10202] = 32'b00000011001001001001100000100000;
   assign mem[10203] = 32'b00000001001000110011000000110100;
   assign mem[10204] = 32'b00000001010111110000100101010110;
   assign mem[10205] = 32'b11111111010100110111010100011001;
   assign mem[10206] = 32'b11110111110101101000110011110000;
   assign mem[10207] = 32'b00000000111001010100001000001011;
   assign mem[10208] = 32'b00000010101011110011101011110100;
   assign mem[10209] = 32'b11110001000000000001001000100000;
   assign mem[10210] = 32'b00000110100110011001011000111000;
   assign mem[10211] = 32'b11110010111111110110101010000000;
   assign mem[10212] = 32'b00000100111100100101100001000000;
   assign mem[10213] = 32'b11110000110111011101010000000000;
   assign mem[10214] = 32'b00000001100001110001100101111010;
   assign mem[10215] = 32'b11111011010111111111001000100000;
   assign mem[10216] = 32'b11111111101010010111100011000011;
   assign mem[10217] = 32'b11111101001010010000111101010100;
   assign mem[10218] = 32'b00000100011101111100110000001000;
   assign mem[10219] = 32'b11111100000101001111100011111100;
   assign mem[10220] = 32'b00000010001001111011001001001100;
   assign mem[10221] = 32'b11111001111110010010110100100000;
   assign mem[10222] = 32'b00000011001100110100001000110100;
   assign mem[10223] = 32'b00000001110110010110010011111000;
   assign mem[10224] = 32'b11111001010111100111010001101000;
   assign mem[10225] = 32'b11111100000101100011010001010100;
   assign mem[10226] = 32'b00000010101000101011101111110100;
   assign mem[10227] = 32'b11111011001001011100011111111000;
   assign mem[10228] = 32'b11111111101101100001000111111110;
   assign mem[10229] = 32'b00000000100011111011011110101011;
   assign mem[10230] = 32'b00000011100110100010110000011100;
   assign mem[10231] = 32'b11111011110111001100101010111000;
   assign mem[10232] = 32'b00000001111010011110011111110000;
   assign mem[10233] = 32'b11110101011110111000110001000000;
   assign mem[10234] = 32'b11111001110100000111111100000000;
   assign mem[10235] = 32'b11111110001001111100000001111010;
   assign mem[10236] = 32'b00000100000101001110100000101000;
   assign mem[10237] = 32'b11111010010110100110100011000000;
   assign mem[10238] = 32'b00000001001010001011110000100100;
   assign mem[10239] = 32'b00000001111110010011011111011100;
   assign mem[10240] = 32'b11111011010000101010011111010000;
   assign mem[10241] = 32'b11111110010010001011000000011000;
   assign mem[10242] = 32'b11111100001001001111011000011100;
   assign mem[10243] = 32'b00000000010010000110100110110001;
   assign mem[10244] = 32'b00000001100000110001101111100100;
   assign mem[10245] = 32'b00000001111000000001110001001110;
   assign mem[10246] = 32'b11111110001101011001110010001100;
   assign mem[10247] = 32'b11111101000001001100001011001000;
   assign mem[10248] = 32'b11111111101111011110010010000011;
   assign mem[10249] = 32'b00000011010010000001111100100100;
   assign mem[10250] = 32'b00000000011111100110110101100100;
   assign mem[10251] = 32'b00000010011011111110111001011000;
   assign mem[10252] = 32'b11100010110000100011011010000000;
   assign mem[10253] = 32'b00001001010101110011111011110000;
   assign mem[10254] = 32'b11111001011000001110110010010000;
   assign mem[10255] = 32'b00000111111010100101010011110000;
   assign mem[10256] = 32'b11101100000000000001111111000000;
   assign mem[10257] = 32'b00001011101010110100110011100000;
   assign mem[10258] = 32'b11100110001110110000001110000000;
   assign mem[10259] = 32'b00000001001001010111011010111110;
   assign mem[10260] = 32'b00000010001110001011101110011000;
   assign mem[10261] = 32'b11110111101101101001101110000000;
   assign mem[10262] = 32'b11111100111010000001001010001100;
   assign mem[10263] = 32'b11111010100000100100001000100000;
   assign mem[10264] = 32'b00000100000110010001110101010000;
   assign mem[10265] = 32'b00000010000100101000010110111100;
   assign mem[10266] = 32'b00000000101101111010011000010010;
   assign mem[10267] = 32'b11110001111000010011110101010000;
   assign mem[10268] = 32'b00000111010101010111101101000000;
   assign mem[10269] = 32'b11111111001110110010001100001000;
   assign mem[10270] = 32'b11110101010101111011101100010000;
   assign mem[10271] = 32'b11110110111110000111101100110000;
   assign mem[10272] = 32'b11110100011011000010001100100000;
   assign mem[10273] = 32'b00000011011010010011110010000000;
   assign mem[10274] = 32'b00000101110011011010110000100000;
   assign mem[10275] = 32'b11111110100000010010001001101000;
   assign mem[10276] = 32'b11101010000100001011111011000000;
   assign mem[10277] = 32'b11111110111101011111101010011010;
   assign mem[10278] = 32'b11111011000011111101111110010000;
   assign mem[10279] = 32'b00000110011000001011000001010000;
   assign mem[10280] = 32'b11101100001001110110111000100000;
   assign mem[10281] = 32'b00000011110000010111111110111000;
   assign mem[10282] = 32'b11111111001001011110000101101111;
   assign mem[10283] = 32'b00000011011011111011110111110000;
   assign mem[10284] = 32'b00000011101110111110110001100000;
   assign mem[10285] = 32'b00000110111111110001010110001000;
   assign mem[10286] = 32'b11011111010000101100100011000000;
   assign mem[10287] = 32'b00000110110100101011110010101000;
   assign mem[10288] = 32'b11111010011111010001010111110000;
   assign mem[10289] = 32'b00000001100000011011001000101010;
   assign mem[10290] = 32'b00000100110111110101111011010000;
   assign mem[10291] = 32'b11111110100000010111110110111000;
   assign mem[10292] = 32'b00000101110110111010011110101000;
   assign mem[10293] = 32'b11110000001101010101001110110000;
   assign mem[10294] = 32'b00000111100100110000100110111000;
   assign mem[10295] = 32'b11111001111000111001110010010000;
   assign mem[10296] = 32'b11111101101110000000011011110100;
   assign mem[10297] = 32'b11111100010001111101110100110000;
   assign mem[10298] = 32'b00000011110010101001011011000000;
   assign mem[10299] = 32'b00000001011100111000011101001000;
   assign mem[10300] = 32'b11111001100101101111111101000000;
   assign mem[10301] = 32'b00001001111110000111000011010000;
   assign mem[10302] = 32'b00000011001001011101110111110100;
   assign mem[10303] = 32'b11111110010001110100101000001110;
   assign mem[10304] = 32'b11110010010010010111000110110000;
   assign mem[10305] = 32'b11111100100001010110001110101100;
   assign mem[10306] = 32'b11111011000000101001000100000000;
   assign mem[10307] = 32'b00001011110111111101010101110000;
   assign mem[10308] = 32'b11111101110000100111101110100000;
   assign mem[10309] = 32'b11110011111110101101010110110000;
   assign mem[10310] = 32'b00000100001110101111001000100000;
   assign mem[10311] = 32'b00000110011000000111100100000000;
   assign mem[10312] = 32'b00000000100011111111011010110110;
   assign mem[10313] = 32'b11111101010011100111110010110100;
   assign mem[10314] = 32'b00000000010100110110110111000001;
   assign mem[10315] = 32'b11111011000100101010001001100000;
   assign mem[10316] = 32'b00000000100100110110010011100011;
   assign mem[10317] = 32'b00001000001001001000110001100000;
   assign mem[10318] = 32'b00001011100001110100101000010000;
   assign mem[10319] = 32'b11100110011110101001010010000000;
   assign mem[10320] = 32'b11101000100110000101001110100000;
   assign mem[10321] = 32'b00000101010110010111001001111000;
   assign mem[10322] = 32'b11111010110101001011011001101000;
   assign mem[10323] = 32'b00001000110100010110101000000000;
   assign mem[10324] = 32'b11111110110000111001001001000000;
   assign mem[10325] = 32'b00000101010010011011000101100000;
   assign mem[10326] = 32'b11100001100001001101011111100000;
   assign mem[10327] = 32'b00000010001000000011100110011100;
   assign mem[10328] = 32'b11110101100111000110111111100000;
   assign mem[10329] = 32'b00000010011100111100010010001000;
   assign mem[10330] = 32'b00000101111100101110100010000000;
   assign mem[10331] = 32'b00000100010001010000111010001000;
   assign mem[10332] = 32'b00000110000000011111000100111000;
   assign mem[10333] = 32'b11110100101111110011000011010000;
   assign mem[10334] = 32'b11111010001010011111010110010000;
   assign mem[10335] = 32'b11111010101110001000100000110000;
   assign mem[10336] = 32'b11111111011010011000100000001011;
   assign mem[10337] = 32'b11111001101001010010110000010000;
   assign mem[10338] = 32'b00000001110000010111011000100110;
   assign mem[10339] = 32'b11111001111100100111000101001000;
   assign mem[10340] = 32'b00000000000000111111011111011101;
   assign mem[10341] = 32'b00001001011010111100001000110000;
   assign mem[10342] = 32'b11111100010011100011111000110000;
   assign mem[10343] = 32'b11111011111011111001000111001000;
   assign mem[10344] = 32'b11111001000000011011001100110000;
   assign mem[10345] = 32'b11111001110011001110011101010000;
   assign mem[10346] = 32'b00000001111001011101011000001100;
   assign mem[10347] = 32'b00000111011100001011000010001000;
   assign mem[10348] = 32'b00000011000100000000001000011000;
   assign mem[10349] = 32'b11111010010100011111111101110000;
   assign mem[10350] = 32'b11111111011010001011011010010001;
   assign mem[10351] = 32'b11110100111000001100011001100000;
   assign mem[10352] = 32'b11110011111100111010011000000000;
   assign mem[10353] = 32'b11111011000011001000000101001000;
   assign mem[10354] = 32'b00000001110110000111011101101000;
   assign mem[10355] = 32'b00000000000110000111000001111000;
   assign mem[10356] = 32'b00000010010101111101001110010000;
   assign mem[10357] = 32'b00000100100011111000110100110000;
   assign mem[10358] = 32'b00000000001010011011000111111101;
   assign mem[10359] = 32'b00001000001000000001100111010000;
   assign mem[10360] = 32'b00000011001100100111101111110000;
   assign mem[10361] = 32'b00000100111100011010011101101000;
   assign mem[10362] = 32'b11111010010110110010010101011000;
   assign mem[10363] = 32'b11110111111110101011010000000000;
   assign mem[10364] = 32'b00000001111010111111000010100000;
   assign mem[10365] = 32'b11111100000001100111100100011000;
   assign mem[10366] = 32'b11111111111111110011111111100100;
   assign mem[10367] = 32'b11111101000110000001101110110000;
   assign mem[10368] = 32'b11111111110000000010011001110110;
   assign mem[10369] = 32'b00001100011110000111011101110000;
   assign mem[10370] = 32'b00000001111010011001000000101000;
   assign mem[10371] = 32'b00001010101101011101100011110000;
   assign mem[10372] = 32'b11111010011100111011001010001000;
   assign mem[10373] = 32'b00000001000100001111000000011010;
   assign mem[10374] = 32'b00000010010111110000111111100000;
   assign mem[10375] = 32'b00000011101110110010010110101100;
   assign mem[10376] = 32'b11111101111101010110001110000000;
   assign mem[10377] = 32'b00000000110001100110010001000110;
   assign mem[10378] = 32'b11111011110100110010010001010000;
   assign mem[10379] = 32'b00000010010010101111000111110100;
   assign mem[10380] = 32'b00000010111110101010011010000000;
   assign mem[10381] = 32'b00000001011001001011000110101100;
   assign mem[10382] = 32'b11111111110000101010101011101010;
   assign mem[10383] = 32'b11111001001110111110001000101000;
   assign mem[10384] = 32'b00000101001100110100010011110000;
   assign mem[10385] = 32'b00000001011101101101001000010010;
   assign mem[10386] = 32'b00000000011011001011110101100001;
   assign mem[10387] = 32'b11110000001100110010101011010000;
   assign mem[10388] = 32'b00000010100110010101110110010100;
   assign mem[10389] = 32'b00000110100101110111000111110000;
   assign mem[10390] = 32'b00000001111101110011001011111010;
   assign mem[10391] = 32'b00000001011110101110111011101110;
   assign mem[10392] = 32'b00000011011101010001011011000000;
   assign mem[10393] = 32'b11111110011101111100011011010010;
   assign mem[10394] = 32'b00000100000110001100010111101000;
   assign mem[10395] = 32'b11111011011010010011110010011000;
   assign mem[10396] = 32'b00000000100010101110100110011111;
   assign mem[10397] = 32'b11111100101011001100100001100000;
   assign mem[10398] = 32'b00000111100011110001011001000000;
   assign mem[10399] = 32'b11111001000000111010111000101000;
   assign mem[10400] = 32'b11111111010001001010101001010111;
   assign mem[10401] = 32'b00000000010111110110010000101101;
   assign mem[10402] = 32'b00000101000101001110000001111000;
   assign mem[10403] = 32'b11111101111011001001100111111000;
   assign mem[10404] = 32'b11111111110010101101101001110001;
   assign mem[10405] = 32'b00000000010010011111110110011101;
   assign mem[10406] = 32'b11111101111010101000101111011100;
   assign mem[10407] = 32'b11111100101011100111011011110000;
   assign mem[10408] = 32'b11110101111111111010110001000000;
   assign mem[10409] = 32'b00000010011100110001000101111100;
   assign mem[10410] = 32'b00000110001101111100100000111000;
   assign mem[10411] = 32'b11111010111101110101011010111000;
   assign mem[10412] = 32'b00000000000110011010100010111011;
   assign mem[10413] = 32'b11110111110101000001010101100000;
   assign mem[10414] = 32'b11111110110101010001101111100000;
   assign mem[10415] = 32'b11110111000101010101100100000000;
   assign mem[10416] = 32'b00000100001100110101011011001000;
   assign mem[10417] = 32'b11111100010010100001011001010100;
   assign mem[10418] = 32'b11111111100100000110010000111100;
   assign mem[10419] = 32'b00000000110001100110110110000010;
   assign mem[10420] = 32'b11111011010100111101000101110000;
   assign mem[10421] = 32'b00000000000000000001001100110110;
   assign mem[10422] = 32'b11111001011100001111100111000000;
   assign mem[10423] = 32'b00000010011000110001001101011100;
   assign mem[10424] = 32'b00001010100011101101000001110000;
   assign mem[10425] = 32'b00000100001000110000101011001000;
   assign mem[10426] = 32'b11110100100110011111000011010000;
   assign mem[10427] = 32'b11111011111000010011101110101000;
   assign mem[10428] = 32'b11111001110001111100110110101000;
   assign mem[10429] = 32'b00000000001000001001001010011101;
   assign mem[10430] = 32'b11111110010101001011001000000010;
   assign mem[10431] = 32'b00000011100011100111111101001000;
   assign mem[10432] = 32'b00000100101110100101111011000000;
   assign mem[10433] = 32'b11111111000110111100110111000000;
   assign mem[10434] = 32'b00000100011111110001001110010000;
   assign mem[10435] = 32'b00000001010001100101010011001000;
   assign mem[10436] = 32'b11110100111000000110101011010000;
   assign mem[10437] = 32'b00000001111110110000111111111010;
   assign mem[10438] = 32'b00000011101001101110011000011100;
   assign mem[10439] = 32'b11111101010111001111101110110100;
   assign mem[10440] = 32'b00000100001000000111001001011000;
   assign mem[10441] = 32'b00000010011010100000100010100000;
   assign mem[10442] = 32'b00000011001100011001010111100100;
   assign mem[10443] = 32'b11110101001001110010010001110000;
   assign mem[10444] = 32'b00000000100100011010001101001100;
   assign mem[10445] = 32'b11111100010001010011010101110100;
   assign mem[10446] = 32'b00000110010011010110010100000000;
   assign mem[10447] = 32'b11111110011001100011011110001000;
   assign mem[10448] = 32'b00000001110000011110010111010100;
   assign mem[10449] = 32'b11111000111100111110111001001000;
   assign mem[10450] = 32'b11111111101101110111011010111110;
   assign mem[10451] = 32'b11111110101101100000100011110000;
   assign mem[10452] = 32'b00000101010011010011111111100000;
   assign mem[10453] = 32'b11111110000001001011011111110010;
   assign mem[10454] = 32'b00000000110110110110010011111100;
   assign mem[10455] = 32'b11111011111011010110110001111000;
   assign mem[10456] = 32'b11111000011111101111010000100000;
   assign mem[10457] = 32'b00000001100010111110011100010100;
   assign mem[10458] = 32'b11111101110011000111000100011000;
   assign mem[10459] = 32'b00000011001011100001010001011100;
   assign mem[10460] = 32'b00000100010011001000001000010000;
   assign mem[10461] = 32'b00000100000001000110100010001000;
   assign mem[10462] = 32'b00000100100110111001110101001000;
   assign mem[10463] = 32'b11110100010010001100101001100000;
   assign mem[10464] = 32'b00000100110011110110111011111000;
   assign mem[10465] = 32'b11111101010111000010001110001100;
   assign mem[10466] = 32'b00000001000001011110110111001000;
   assign mem[10467] = 32'b11110110110100111011001111110000;
   assign mem[10468] = 32'b00001000100011100001110001110000;
   assign mem[10469] = 32'b11111000110010101000011101100000;
   assign mem[10470] = 32'b00000100011110111011001011110000;
   assign mem[10471] = 32'b11110100011100110110011010010000;
   assign mem[10472] = 32'b00000010111110011101011010111100;
   assign mem[10473] = 32'b11111111111100010110010101101101;
   assign mem[10474] = 32'b00000001111101101100010110010110;
   assign mem[10475] = 32'b11111011001110110110110001000000;
   assign mem[10476] = 32'b00000101000100111111101101011000;
   assign mem[10477] = 32'b11111011000101000000011000001000;
   assign mem[10478] = 32'b00000001111100001101111101010000;
   assign mem[10479] = 32'b11111111110100111111000000110101;
   assign mem[10480] = 32'b00000001100011100010011001000110;
   assign mem[10481] = 32'b11110011000011011110001011110000;
   assign mem[10482] = 32'b11111111111010011110001001110101;
   assign mem[10483] = 32'b11111001111100000110001010010000;
   assign mem[10484] = 32'b11111110001111001110000111001100;
   assign mem[10485] = 32'b00000001001100011111101101101000;
   assign mem[10486] = 32'b11111110001101110010101001000100;
   assign mem[10487] = 32'b11111001100100110110100111111000;
   assign mem[10488] = 32'b00000110000001111011111001111000;
   assign mem[10489] = 32'b00000100001101101110110100111000;
   assign mem[10490] = 32'b00000100011011110001101101101000;
   assign mem[10491] = 32'b11111101000111111001010001000000;
   assign mem[10492] = 32'b11110111100111000111100110100000;
   assign mem[10493] = 32'b11110101101001011000011010000000;
   assign mem[10494] = 32'b00000111001111100111101011101000;
   assign mem[10495] = 32'b11111000110111111100000000100000;
   assign mem[10496] = 32'b11111011001111000101001011100000;
   assign mem[10497] = 32'b00010011000001110001101001000000;
   assign mem[10498] = 32'b11111111011111010010011100010001;
   assign mem[10499] = 32'b11110111010011110110110100000000;
   assign mem[10500] = 32'b00000010110101011000000101111000;
   assign mem[10501] = 32'b00000100000001101011110001110000;
   assign mem[10502] = 32'b11111001010100000011110111111000;
   assign mem[10503] = 32'b11110111111110011110100010110000;
   assign mem[10504] = 32'b11111110110011011101100111111000;
   assign mem[10505] = 32'b11110101001100100001110101000000;
   assign mem[10506] = 32'b00000101010110111101011000000000;
   assign mem[10507] = 32'b00000100000000010011110001010000;
   assign mem[10508] = 32'b00000001000101101000110010110100;
   assign mem[10509] = 32'b00000111111011101010011001000000;
   assign mem[10510] = 32'b11111001001011001011001110010000;
   assign mem[10511] = 32'b00000011100110101100101000110000;
   assign mem[10512] = 32'b00000111000010000110110000011000;
   assign mem[10513] = 32'b11111111001000000100011000010000;
   assign mem[10514] = 32'b11111001010111001000000011011000;
   assign mem[10515] = 32'b11110110011100110001000111110000;
   assign mem[10516] = 32'b11110100111010001101110100110000;
   assign mem[10517] = 32'b00000110100101101110010100000000;
   assign mem[10518] = 32'b00001000000100111101011001000000;
   assign mem[10519] = 32'b00000000111111011100001111101111;
   assign mem[10520] = 32'b00000010100001101010111101000100;
   assign mem[10521] = 32'b00000010110111011001101011100000;
   assign mem[10522] = 32'b00000011011011001110100111100100;
   assign mem[10523] = 32'b11111000100000101110111010110000;
   assign mem[10524] = 32'b00000010010101000101101101110000;
   assign mem[10525] = 32'b11111100100010101010001011000100;
   assign mem[10526] = 32'b11110111011110100011000101010000;
   assign mem[10527] = 32'b11110101000100101100111110100000;
   assign mem[10528] = 32'b00000001000010000110111111010100;
   assign mem[10529] = 32'b00001000000011111110010010000000;
   assign mem[10530] = 32'b11110010011101111000101011110000;
   assign mem[10531] = 32'b00001000001011010000001011110000;
   assign mem[10532] = 32'b00000001001001000111011010100110;
   assign mem[10533] = 32'b00000011010100111100100001100000;
   assign mem[10534] = 32'b11110011111101011110010011110000;
   assign mem[10535] = 32'b00001000101001110000101100110000;
   assign mem[10536] = 32'b11111001101001001011001011010000;
   assign mem[10537] = 32'b00000110110011000100101010010000;
   assign mem[10538] = 32'b11110011010100110001000000010000;
   assign mem[10539] = 32'b00000000111100101010010101011100;
   assign mem[10540] = 32'b00000000010000110101000000110000;
   assign mem[10541] = 32'b00000000101001000001001110110111;
   assign mem[10542] = 32'b11111101010010000111110110111000;
   assign mem[10543] = 32'b00000001011101010100100100001100;
   assign mem[10544] = 32'b00000101100110100101000011001000;
   assign mem[10545] = 32'b11111011110001000100001011010000;
   assign mem[10546] = 32'b00000010101101001010011110011000;
   assign mem[10547] = 32'b00000000011000000100100111110111;
   assign mem[10548] = 32'b11111010110011110011000101100000;
   assign mem[10549] = 32'b11111110111010100011111000001110;
   assign mem[10550] = 32'b00000001000100000000110101101010;
   assign mem[10551] = 32'b11110111100101001000111100100000;
   assign mem[10552] = 32'b11111011010001101111011010111000;
   assign mem[10553] = 32'b11111100011100010110110011111000;
   assign mem[10554] = 32'b00000100001010100110110011010000;
   assign mem[10555] = 32'b00000010110110011001110100001000;
   assign mem[10556] = 32'b11111001101101110000111001000000;
   assign mem[10557] = 32'b00000001011001001111010000000010;
   assign mem[10558] = 32'b11111011101011100011011111001000;
   assign mem[10559] = 32'b00000011101010011111110110101100;
   assign mem[10560] = 32'b00000110011001100010000100111000;
   assign mem[10561] = 32'b00000101001000110101101101111000;
   assign mem[10562] = 32'b00001000110010101000011010100000;
   assign mem[10563] = 32'b11110011111110000100001110010000;
   assign mem[10564] = 32'b11111101111010110001111011001000;
   assign mem[10565] = 32'b11110101000000111000000011110000;
   assign mem[10566] = 32'b11111111000010000000010110000100;
   assign mem[10567] = 32'b00000000011010100110011000100110;
   assign mem[10568] = 32'b00001011100001011110101001000000;
   assign mem[10569] = 32'b11100111101011010011110001100000;
   assign mem[10570] = 32'b00000100100110110100110001001000;
   assign mem[10571] = 32'b11111101100110000101000001101000;
   assign mem[10572] = 32'b00000100110100000010110011010000;
   assign mem[10573] = 32'b11110100001101100001111010000000;
   assign mem[10574] = 32'b00000110101100001010111001010000;
   assign mem[10575] = 32'b11110110100001110111110100110000;
   assign mem[10576] = 32'b00000111001011100010010100001000;
   assign mem[10577] = 32'b11111100010100101000101111110100;
   assign mem[10578] = 32'b00000100111110111100100111110000;
   assign mem[10579] = 32'b00000001101110111000001101100110;
   assign mem[10580] = 32'b00000010110101001010110100010000;
   assign mem[10581] = 32'b11111101101111010110101010000100;
   assign mem[10582] = 32'b11111101111011100001001111010100;
   assign mem[10583] = 32'b11110110011000011111110011000000;
   assign mem[10584] = 32'b00000100010000110011011000010000;
   assign mem[10585] = 32'b11111100000010111000110101001000;
   assign mem[10586] = 32'b11111000110110110000101111101000;
   assign mem[10587] = 32'b11111110001000111010101111000110;
   assign mem[10588] = 32'b11111110110110000000001000111000;
   assign mem[10589] = 32'b00001000011001001101101000010000;
   assign mem[10590] = 32'b11111001101110011000001100101000;
   assign mem[10591] = 32'b11111111101001010101101000100111;
   assign mem[10592] = 32'b00000101110000011111101110110000;
   assign mem[10593] = 32'b11111011011100010001011110100000;
   assign mem[10594] = 32'b11111000000010100111001111001000;
   assign mem[10595] = 32'b11111001000011111101000100110000;
   assign mem[10596] = 32'b11111100010001100101011010010100;
   assign mem[10597] = 32'b00001011101110111111010000000000;
   assign mem[10598] = 32'b00000010100110001111100010111000;
   assign mem[10599] = 32'b11111000011011100000110000110000;
   assign mem[10600] = 32'b11111101001011100111111000111000;
   assign mem[10601] = 32'b00000011000000001001010011110100;
   assign mem[10602] = 32'b11111000100100101110011101110000;
   assign mem[10603] = 32'b00000101101010110101000111111000;
   assign mem[10604] = 32'b00000110011111100011100000111000;
   assign mem[10605] = 32'b00000101010001000000110000110000;
   assign mem[10606] = 32'b11110101001001010010000100100000;
   assign mem[10607] = 32'b00000000010101010111101110000100;
   assign mem[10608] = 32'b11110111010000011011111101000000;
   assign mem[10609] = 32'b11111111101100101011100110111101;
   assign mem[10610] = 32'b11111101010010101000100011011100;
   assign mem[10611] = 32'b11111110110011001101010000010000;
   assign mem[10612] = 32'b11111100010101101000100100010100;
   assign mem[10613] = 32'b00001000001000100001010111110000;
   assign mem[10614] = 32'b11111111000110000110001011111010;
   assign mem[10615] = 32'b00000101010101010101000101101000;
   assign mem[10616] = 32'b11111110001100101111110111001110;
   assign mem[10617] = 32'b00000101111000011101101011011000;
   assign mem[10618] = 32'b11101110110100010000100110100000;
   assign mem[10619] = 32'b00000011010111100110000000110100;
   assign mem[10620] = 32'b11111101111010111110001010010100;
   assign mem[10621] = 32'b11111100011111110111010110101100;
   assign mem[10622] = 32'b00000001010000001101011111111110;
   assign mem[10623] = 32'b11111001100101001011011111111000;
   assign mem[10624] = 32'b00000011000010011110100100001000;
   assign mem[10625] = 32'b00000010110000111101111111111100;
   assign mem[10626] = 32'b00000010010111000000011000011000;
   assign mem[10627] = 32'b11110010110111001000111101100000;
   assign mem[10628] = 32'b00000000001100000001000000111000;
   assign mem[10629] = 32'b00000111100010011001010111001000;
   assign mem[10630] = 32'b11100100011001101000100001000000;
   assign mem[10631] = 32'b00001000000001111001110000010000;
   assign mem[10632] = 32'b11111110111100011101110011011010;
   assign mem[10633] = 32'b00000000111001100000110010001111;
   assign mem[10634] = 32'b00000011010010011101001010101100;
   assign mem[10635] = 32'b00000110011111111010101111001000;
   assign mem[10636] = 32'b11011111111100000100101100000000;
   assign mem[10637] = 32'b00000011110110111100110010000100;
   assign mem[10638] = 32'b11111000101111010001011011010000;
   assign mem[10639] = 32'b00000001111000000000010100010100;
   assign mem[10640] = 32'b00000101010011011000110110100000;
   assign mem[10641] = 32'b11101110111001010010011011100000;
   assign mem[10642] = 32'b00000001000010010010000100011110;
   assign mem[10643] = 32'b11101111100100100011001110100000;
   assign mem[10644] = 32'b00000011011101001001101100110000;
   assign mem[10645] = 32'b11111100011110010010111011011000;
   assign mem[10646] = 32'b00000101001011000001010010101000;
   assign mem[10647] = 32'b11111100010010100110011101000100;
   assign mem[10648] = 32'b00000001000101001111111110101010;
   assign mem[10649] = 32'b00000110001110110110111010111000;
   assign mem[10650] = 32'b11111011110010110010010000010000;
   assign mem[10651] = 32'b00000000110011110110001110110110;
   assign mem[10652] = 32'b00000101110100111111100001010000;
   assign mem[10653] = 32'b00000010000100010011000010010100;
   assign mem[10654] = 32'b00000010101010111011000000111100;
   assign mem[10655] = 32'b00000101010000011001000100000000;
   assign mem[10656] = 32'b11110111110000111110000000010000;
   assign mem[10657] = 32'b00000011000100010110100001011100;
   assign mem[10658] = 32'b11111100100001001010001001010100;
   assign mem[10659] = 32'b00000011001100001010111111000100;
   assign mem[10660] = 32'b11111001110000101000101100011000;
   assign mem[10661] = 32'b00000001010010110100101101110010;
   assign mem[10662] = 32'b11111001100110110011001100101000;
   assign mem[10663] = 32'b00000110111011110101111011111000;
   assign mem[10664] = 32'b00000100000010011011010100001000;
   assign mem[10665] = 32'b00000011100001110111000101011000;
   assign mem[10666] = 32'b11110100001001111100000010110000;
   assign mem[10667] = 32'b00000100000111101100000110010000;
   assign mem[10668] = 32'b11110111001101100111101110100000;
   assign mem[10669] = 32'b00000101011111100100001101110000;
   assign mem[10670] = 32'b00000000011011101111101100001010;
   assign mem[10671] = 32'b11110100101111100011100001000000;
   assign mem[10672] = 32'b11110100010010101010000010010000;
   assign mem[10673] = 32'b00001101101010110111110101010000;
   assign mem[10674] = 32'b00000000111110000001000010011001;
   assign mem[10675] = 32'b00001000001010010101110000000000;
   assign mem[10676] = 32'b00000010111011100100100010100000;
   assign mem[10677] = 32'b00000001010010010101010011010110;
   assign mem[10678] = 32'b11110100000010101110000000010000;
   assign mem[10679] = 32'b00000001110010011001101110100110;
   assign mem[10680] = 32'b00000001110011111000000100110010;
   assign mem[10681] = 32'b11110100111000100111101110100000;
   assign mem[10682] = 32'b00000011001101100000111010001000;
   assign mem[10683] = 32'b11111011100010111001110100001000;
   assign mem[10684] = 32'b00000100111110011100010111010000;
   assign mem[10685] = 32'b11111110100100000101100110011010;
   assign mem[10686] = 32'b11111110111110110000000110010010;
   assign mem[10687] = 32'b11110011101111110111000110110000;
   assign mem[10688] = 32'b00000011111110000100111101111100;
   assign mem[10689] = 32'b00000001011011001000111111110000;
   assign mem[10690] = 32'b00000000101110010000111110011110;
   assign mem[10691] = 32'b11111000011111111001010000001000;
   assign mem[10692] = 32'b11110011100001110011000000100000;
   assign mem[10693] = 32'b00001000111001100001010101100000;
   assign mem[10694] = 32'b11110110100001011011011111100000;
   assign mem[10695] = 32'b11111001001101100100011011011000;
   assign mem[10696] = 32'b00000100111100000100001111101000;
   assign mem[10697] = 32'b11111101001100110111111000100000;
   assign mem[10698] = 32'b00000100011001000000100000010000;
   assign mem[10699] = 32'b00000001001011000110011100111000;
   assign mem[10700] = 32'b00000101110101111101011110101000;
   assign mem[10701] = 32'b00000011110001010101001011101100;
   assign mem[10702] = 32'b11110101100101011001010011010000;
   assign mem[10703] = 32'b11111000011111101010010111111000;
   assign mem[10704] = 32'b00000100110100111010001111110000;
   assign mem[10705] = 32'b11111000101101011001110111010000;
   assign mem[10706] = 32'b00000011011010101101000101010100;
   assign mem[10707] = 32'b11111010001111011000010101110000;
   assign mem[10708] = 32'b00001001110010000100010010100000;
   assign mem[10709] = 32'b11111111011101010110000101110001;
   assign mem[10710] = 32'b00000010011010100111110000001100;
   assign mem[10711] = 32'b00000001100101100101010010010010;
   assign mem[10712] = 32'b11111110000001001111011010010100;
   assign mem[10713] = 32'b00000011010111100000101111100100;
   assign mem[10714] = 32'b11111101111100110110100011101000;
   assign mem[10715] = 32'b00000011001110101001011010010000;
   assign mem[10716] = 32'b00000011001010101110010110010000;
   assign mem[10717] = 32'b00000010011010100010100001101100;
   assign mem[10718] = 32'b00000011000101001101011010001100;
   assign mem[10719] = 32'b00000000011001001110001110011100;
   assign mem[10720] = 32'b00000001000001110000010000110100;
   assign mem[10721] = 32'b11111001010101111000010000111000;
   assign mem[10722] = 32'b00000110010101111001110011011000;
   assign mem[10723] = 32'b11111101110110110000101101000100;
   assign mem[10724] = 32'b00000100000010011101110001011000;
   assign mem[10725] = 32'b11111001000110001011001101110000;
   assign mem[10726] = 32'b00000011001110001110000100100000;
   assign mem[10727] = 32'b11111100001010111001101101010100;
   assign mem[10728] = 32'b00000101110110100011101001101000;
   assign mem[10729] = 32'b11111111111011100000100110000001;
   assign mem[10730] = 32'b11111111000111101001010111001100;
   assign mem[10731] = 32'b00000100010001001001111110011000;
   assign mem[10732] = 32'b00000110000001000011101111110000;
   assign mem[10733] = 32'b11110100010100100100100000010000;
   assign mem[10734] = 32'b11110111110111011100101010000000;
   assign mem[10735] = 32'b11110011110100000001000111110000;
   assign mem[10736] = 32'b11111111011110001000000001101100;
   assign mem[10737] = 32'b00000000011010001000101110010110;
   assign mem[10738] = 32'b00001000010101100010111000010000;
   assign mem[10739] = 32'b11111011100111000100010010011000;
   assign mem[10740] = 32'b00000000001001001100000001011010;
   assign mem[10741] = 32'b11111000001110001111101000010000;
   assign mem[10742] = 32'b00000101110010011100010011001000;
   assign mem[10743] = 32'b11110000001101110010101001000000;
   assign mem[10744] = 32'b00000011001111101001011100011100;
   assign mem[10745] = 32'b11111011111001011101110111000000;
   assign mem[10746] = 32'b11111000000010111100000111010000;
   assign mem[10747] = 32'b00000010101011111110101000010100;
   assign mem[10748] = 32'b00001001100110110001100111110000;
   assign mem[10749] = 32'b11111010000001010000001011000000;
   assign mem[10750] = 32'b00000011011110101011000001100100;
   assign mem[10751] = 32'b00000001011111000011110100000010;
   assign mem[10752] = 32'b11111100110000101000101000100000;
   assign mem[10753] = 32'b00001111011110110010100000100000;
   assign mem[10754] = 32'b11111010000011100001011101011000;
   assign mem[10755] = 32'b00000100001111110001010101110000;
   assign mem[10756] = 32'b11111110010001000111101001101010;
   assign mem[10757] = 32'b11111010110111000010011110101000;
   assign mem[10758] = 32'b00000000010000001011101001011111;
   assign mem[10759] = 32'b11111111101010011011100000010111;
   assign mem[10760] = 32'b11111110010110010001011000011010;
   assign mem[10761] = 32'b11111111011101110000010010011000;
   assign mem[10762] = 32'b00000000011010001010000011010000;
   assign mem[10763] = 32'b11111111110010001111000001110111;
   assign mem[10764] = 32'b00000001011101111110100001000010;
   assign mem[10765] = 32'b11111111100100100010110101011011;
   assign mem[10766] = 32'b11111101110010001001000101111000;
   assign mem[10767] = 32'b11111100011001000100111110101000;
   assign mem[10768] = 32'b11111011101100000101000001101000;
   assign mem[10769] = 32'b00000011001111010100100101011100;
   assign mem[10770] = 32'b00000000100111001011101111111110;
   assign mem[10771] = 32'b00000010100101110001010100010100;
   assign mem[10772] = 32'b11111110101010111111110011001110;
   assign mem[10773] = 32'b11111100110111111110101001001000;
   assign mem[10774] = 32'b00001011000010011000100010000000;
   assign mem[10775] = 32'b11111110011100100111100100001100;
   assign mem[10776] = 32'b11111001110010110010001010010000;
   assign mem[10777] = 32'b00000010111110010111000011010000;
   assign mem[10778] = 32'b11111011001000010010010001100000;
   assign mem[10779] = 32'b00000100001110100110110111100000;
   assign mem[10780] = 32'b11111111111010111110011100111111;
   assign mem[10781] = 32'b11111110011100100101110110011000;
   assign mem[10782] = 32'b00000001001000001010111100011010;
   assign mem[10783] = 32'b11111010110001011100100011001000;
   assign mem[10784] = 32'b00000100001010001000100100010000;
   assign mem[10785] = 32'b00000011000110000110010101010100;
   assign mem[10786] = 32'b11111110101111110010001010101110;
   assign mem[10787] = 32'b00000001110110111010100110111000;
   assign mem[10788] = 32'b11111100010001110110011011110100;
   assign mem[10789] = 32'b00000000111110101000100111111110;
   assign mem[10790] = 32'b00000111001101111110001100000000;
   assign mem[10791] = 32'b00000011110111000001010001110100;
   assign mem[10792] = 32'b11111010110100101110111001111000;
   assign mem[10793] = 32'b11110111000110010110110110100000;
   assign mem[10794] = 32'b11111011000111000010010111010000;
   assign mem[10795] = 32'b11111010011010101011010001111000;
   assign mem[10796] = 32'b00000110011000010011100101111000;
   assign mem[10797] = 32'b11111110100001111101101010101100;
   assign mem[10798] = 32'b00000000011010111101011110011101;
   assign mem[10799] = 32'b11111011001101000101111010001000;
   assign mem[10800] = 32'b11111110111100000001001100010100;
   assign mem[10801] = 32'b11111010101010110100101101110000;
   assign mem[10802] = 32'b00000110000101101001000111100000;
   assign mem[10803] = 32'b00000010001011110001100011100100;
   assign mem[10804] = 32'b11111111101110011011011101101100;
   assign mem[10805] = 32'b11111110010101101111011000010110;
   assign mem[10806] = 32'b11111101011101001011101000010100;
   assign mem[10807] = 32'b00000100110110110111010101111000;
   assign mem[10808] = 32'b00000011101011001110111010111000;
   assign mem[10809] = 32'b11111001101011100111100100111000;
   assign mem[10810] = 32'b11111010110011101111011010010000;
   assign mem[10811] = 32'b11110000111000010011100101010000;
   assign mem[10812] = 32'b11110000010000000110010101110000;
   assign mem[10813] = 32'b11111101011000011010011011110000;
   assign mem[10814] = 32'b00000100101011000001101010011000;
   assign mem[10815] = 32'b00000001000110000101011101000010;
   assign mem[10816] = 32'b11111111101111011110101011110101;
   assign mem[10817] = 32'b11111101001011000111101110011000;
   assign mem[10818] = 32'b00000011110110100001100010111100;
   assign mem[10819] = 32'b00000110001010110001111011110000;
   assign mem[10820] = 32'b11111111011111111100100110010100;
   assign mem[10821] = 32'b00000101000001001000111000011000;
   assign mem[10822] = 32'b00000000111001000101011000101000;
   assign mem[10823] = 32'b00001000010010011001001011010000;
   assign mem[10824] = 32'b11111010010000011101011010001000;
   assign mem[10825] = 32'b00001001111100011001100011110000;
   assign mem[10826] = 32'b11110110010000100101011000110000;
   assign mem[10827] = 32'b00000010010011010001001000010100;
   assign mem[10828] = 32'b11101110001001111101010101000000;
   assign mem[10829] = 32'b11111110110111001111001101010110;
   assign mem[10830] = 32'b11111101101101000111111010000100;
   assign mem[10831] = 32'b00000001001001001000000000101100;
   assign mem[10832] = 32'b00000001010000100100111000101000;
   assign mem[10833] = 32'b00001010010100000110000110100000;
   assign mem[10834] = 32'b11110111110101011001100011110000;
   assign mem[10835] = 32'b00000011101101111011011000000100;
   assign mem[10836] = 32'b11111111101011011101110110110000;
   assign mem[10837] = 32'b11111100101110111111011001110000;
   assign mem[10838] = 32'b00000001000011110011101100011010;
   assign mem[10839] = 32'b11111100110011100000111110100100;
   assign mem[10840] = 32'b11110011101010101101001010000000;
   assign mem[10841] = 32'b11111111110110001101010111110110;
   assign mem[10842] = 32'b00000011101010010000001000100000;
   assign mem[10843] = 32'b11111111001001101111000100001100;
   assign mem[10844] = 32'b11111100011011111110111111110000;
   assign mem[10845] = 32'b00000010001110000100101101100000;
   assign mem[10846] = 32'b11101111001010100101110110100000;
   assign mem[10847] = 32'b00000101101001101001010010001000;
   assign mem[10848] = 32'b11111101010110110000000011000100;
   assign mem[10849] = 32'b00000000000110100011011100111010;
   assign mem[10850] = 32'b00000110001001000010110111011000;
   assign mem[10851] = 32'b00000011001011010000111101010100;
   assign mem[10852] = 32'b00001000001001001110000010110000;
   assign mem[10853] = 32'b11111010100011010000101101101000;
   assign mem[10854] = 32'b11111001011100011001001101000000;
   assign mem[10855] = 32'b11110100000010011000100000010000;
   assign mem[10856] = 32'b00000001010111010001100001100000;
   assign mem[10857] = 32'b00000000110001101011001110101001;
   assign mem[10858] = 32'b00001000011100101001101001100000;
   assign mem[10859] = 32'b11111101011101110001110100010100;
   assign mem[10860] = 32'b00000100000010011000111110000000;
   assign mem[10861] = 32'b11111111001010110101101110011110;
   assign mem[10862] = 32'b00000101111111110100101011101000;
   assign mem[10863] = 32'b11111101101100100011110101000100;
   assign mem[10864] = 32'b00000000001010111011101001010001;
   assign mem[10865] = 32'b11111101000100011011000001101100;
   assign mem[10866] = 32'b00000011011001000111110100011000;
   assign mem[10867] = 32'b11110110000100010011010010110000;
   assign mem[10868] = 32'b11111111011100101011101001111110;
   assign mem[10869] = 32'b00000010110010011011110000000000;
   assign mem[10870] = 32'b00000100000000111101011100100000;
   assign mem[10871] = 32'b00000010111101110010011100011100;
   assign mem[10872] = 32'b00000111100100100010101110010000;
   assign mem[10873] = 32'b11110100101010000011101100010000;
   assign mem[10874] = 32'b00000001001010010010101011100110;
   assign mem[10875] = 32'b11111100000001000100000011010000;
   assign mem[10876] = 32'b00000010101101011000011000111100;
   assign mem[10877] = 32'b11111010101111011000000001000000;
   assign mem[10878] = 32'b00001000000110111110110100000000;
   assign mem[10879] = 32'b11111011001011111000011000000000;
   assign mem[10880] = 32'b11111010110001000100000001101000;
   assign mem[10881] = 32'b00000000100001010010010001011001;
   assign mem[10882] = 32'b00000100010001001101101010001000;
   assign mem[10883] = 32'b00000111011001100111110011011000;
   assign mem[10884] = 32'b11111111000010011101000011111100;
   assign mem[10885] = 32'b00000011000010101001000110101100;
   assign mem[10886] = 32'b11111111010110111001100000101011;
   assign mem[10887] = 32'b11110010100110010111010101100000;
   assign mem[10888] = 32'b00000100001111101001101110010000;
   assign mem[10889] = 32'b11111111011000101100101010001110;
   assign mem[10890] = 32'b00010001000111011100111110100000;
   assign mem[10891] = 32'b00000101001110100111000101110000;
   assign mem[10892] = 32'b11101011110011011010110111000000;
   assign mem[10893] = 32'b00001000010010000100010010100000;
   assign mem[10894] = 32'b11111010100010101011111001010000;
   assign mem[10895] = 32'b00001010110001100100010001010000;
   assign mem[10896] = 32'b11111001010101110010000001000000;
   assign mem[10897] = 32'b00001111100110101011001110100000;
   assign mem[10898] = 32'b11100011111111010010001101100000;
   assign mem[10899] = 32'b11111000110110101000001011000000;
   assign mem[10900] = 32'b11111110100010010100110101000010;
   assign mem[10901] = 32'b11110000001100010100100010100000;
   assign mem[10902] = 32'b00000100001101111000001111100000;
   assign mem[10903] = 32'b00000000111111100101011001001111;
   assign mem[10904] = 32'b00000011001001101111010010010100;
   assign mem[10905] = 32'b00000001010011100110010011111010;
   assign mem[10906] = 32'b00000001110000110100010010011000;
   assign mem[10907] = 32'b11101101000111100001010101000000;
   assign mem[10908] = 32'b00000010101101110010111011011000;
   assign mem[10909] = 32'b00000000111101110011110010011010;
   assign mem[10910] = 32'b11110011001011100011000110010000;
   assign mem[10911] = 32'b11100110101010101100010110000000;
   assign mem[10912] = 32'b00000001010110111110010011001100;
   assign mem[10913] = 32'b00000000010001001001110100011000;
   assign mem[10914] = 32'b00000111100111111101000010100000;
   assign mem[10915] = 32'b00000000100110010110010101001110;
   assign mem[10916] = 32'b11110011001000100101100000010000;
   assign mem[10917] = 32'b11111011010010101111100000101000;
   assign mem[10918] = 32'b11111011010110010011011000011000;
   assign mem[10919] = 32'b00001010111010111011010101000000;
   assign mem[10920] = 32'b11110101011001001011010000100000;
   assign mem[10921] = 32'b11111101101010000110001110101100;
   assign mem[10922] = 32'b11111100110010110111110101110100;
   assign mem[10923] = 32'b00000010000011101001111010101100;
   assign mem[10924] = 32'b00000101111010001010111110001000;
   assign mem[10925] = 32'b00000000010100100000010111101011;
   assign mem[10926] = 32'b11110011110010001001110110010000;
   assign mem[10927] = 32'b11111010011111001110000000010000;
   assign mem[10928] = 32'b11111001001011000110100111101000;
   assign mem[10929] = 32'b00000111000101101110101111111000;
   assign mem[10930] = 32'b00000001010010001110001000111010;
   assign mem[10931] = 32'b00000010011111001001111000010100;
   assign mem[10932] = 32'b00000000000001000011101100001011;
   assign mem[10933] = 32'b11111010101111110111100011110000;
   assign mem[10934] = 32'b00000111001100011011001101100000;
   assign mem[10935] = 32'b11110111011001110101101000010000;
   assign mem[10936] = 32'b00000100111010011100011100011000;
   assign mem[10937] = 32'b11111100101000011011001011111100;
   assign mem[10938] = 32'b00000100100110110101110010111000;
   assign mem[10939] = 32'b11111101010010010001111001111100;
   assign mem[10940] = 32'b00000101100011111011011011110000;
   assign mem[10941] = 32'b00010000111100100100010100000000;
   assign mem[10942] = 32'b11111100101111100101010111111000;
   assign mem[10943] = 32'b11110110111011001010100011010000;
   assign mem[10944] = 32'b11110111111000111001110100000000;
   assign mem[10945] = 32'b00000001111010001011110111100100;
   assign mem[10946] = 32'b11110110111101101101110111010000;
   assign mem[10947] = 32'b00001100110010001000111011010000;
   assign mem[10948] = 32'b11111100100001011011011110111100;
   assign mem[10949] = 32'b11110111001010111001111110010000;
   assign mem[10950] = 32'b00000000011101010011000011010011;
   assign mem[10951] = 32'b00000000101110101101101011000010;
   assign mem[10952] = 32'b00000011100011110011000010000100;
   assign mem[10953] = 32'b11111110011101001011101100101000;
   assign mem[10954] = 32'b11111011010010011010010010010000;
   assign mem[10955] = 32'b11111100011011000100100100110100;
   assign mem[10956] = 32'b11111000011111101011001010101000;
   assign mem[10957] = 32'b11111111001101011100101001010110;
   assign mem[10958] = 32'b11111111000001010010011111011111;
   assign mem[10959] = 32'b00001000110001101110111110010000;
   assign mem[10960] = 32'b00000001001110111011101011101110;
   assign mem[10961] = 32'b00001011100000001100010010000000;
   assign mem[10962] = 32'b11111000011011101101110000010000;
   assign mem[10963] = 32'b00001000010011111011001111010000;
   assign mem[10964] = 32'b11111011100011010001111100101000;
   assign mem[10965] = 32'b11111110111111110100111101110000;
   assign mem[10966] = 32'b11110101011111100010010100000000;
   assign mem[10967] = 32'b00000100010011100001110101110000;
   assign mem[10968] = 32'b11101001010000110110011110100000;
   assign mem[10969] = 32'b11111110101000110110101001000110;
   assign mem[10970] = 32'b00000100011011100000110001101000;
   assign mem[10971] = 32'b00000100011100000010110100110000;
   assign mem[10972] = 32'b11111100110010011100001100110000;
   assign mem[10973] = 32'b11111010110111000001101010101000;
   assign mem[10974] = 32'b11111111011100110001101100001001;
   assign mem[10975] = 32'b00000010110000100011000101101000;
   assign mem[10976] = 32'b11111000110000001111010011111000;
   assign mem[10977] = 32'b00000011111001000111111100010000;
   assign mem[10978] = 32'b11111011100110101111011101011000;
   assign mem[10979] = 32'b00000000110011111010100001001011;
   assign mem[10980] = 32'b11111100110110110110001010011000;
   assign mem[10981] = 32'b00000000101011100001111001110010;
   assign mem[10982] = 32'b11111101100101000000010101111000;
   assign mem[10983] = 32'b11111101011011000111100000000000;
   assign mem[10984] = 32'b00000100101110000011110110101000;
   assign mem[10985] = 32'b00000000000100010011001100010010;
   assign mem[10986] = 32'b11111010000111011100001010100000;
   assign mem[10987] = 32'b11111101010111100110010100100100;
   assign mem[10988] = 32'b00000001100011000011110000110010;
   assign mem[10989] = 32'b00000111001110100110111100011000;
   assign mem[10990] = 32'b00000010101100101100111101000100;
   assign mem[10991] = 32'b00000101111001001100001110000000;
   assign mem[10992] = 32'b00000000010011111000001101011000;
   assign mem[10993] = 32'b00000111101001100001100000011000;
   assign mem[10994] = 32'b11111101111000101010011001011000;
   assign mem[10995] = 32'b00000001001011101010010100011100;
   assign mem[10996] = 32'b11111101011011010111111101001000;
   assign mem[10997] = 32'b11111101001001000111111110000000;
   assign mem[10998] = 32'b11111101011100010011001101100100;
   assign mem[10999] = 32'b11111110000001011010100000111110;
   assign mem[11000] = 32'b00000001001010100100001100001000;
   assign mem[11001] = 32'b00000011011101000001111111001100;
   assign mem[11002] = 32'b11111100000100001011110111011100;
   assign mem[11003] = 32'b11110110000100110011100001110000;
   assign mem[11004] = 32'b00001101000001110011001001000000;
   assign mem[11005] = 32'b11111100100100010100101011010100;
   assign mem[11006] = 32'b00000010010111011110010110111100;
   assign mem[11007] = 32'b11110111001010000000110000110000;
   assign mem[11008] = 32'b11111000110011011111101011101000;
   assign mem[11009] = 32'b00001101000010100111101101110000;
   assign mem[11010] = 32'b11111110011001100100000110000110;
   assign mem[11011] = 32'b11111111110100111001101111001000;
   assign mem[11012] = 32'b11111111000011010101101011010100;
   assign mem[11013] = 32'b00000001000101101010100110100000;
   assign mem[11014] = 32'b00000110010101000101010101101000;
   assign mem[11015] = 32'b11111111100011111100111111000110;
   assign mem[11016] = 32'b00000110010010110000000001110000;
   assign mem[11017] = 32'b11110110010100110101110010000000;
   assign mem[11018] = 32'b11111001100111111110100100010000;
   assign mem[11019] = 32'b11111101111101010111011101111000;
   assign mem[11020] = 32'b00000010100100101101000010000100;
   assign mem[11021] = 32'b11110111000110100100101100000000;
   assign mem[11022] = 32'b00000110011010001101000100000000;
   assign mem[11023] = 32'b11111110110011111100001010001100;
   assign mem[11024] = 32'b00000101000000100110010111100000;
   assign mem[11025] = 32'b11111010101010000010100000010000;
   assign mem[11026] = 32'b00000001011111001000001000101000;
   assign mem[11027] = 32'b11110001001101010010101000100000;
   assign mem[11028] = 32'b00000000010001110110001100001010;
   assign mem[11029] = 32'b00000010101110101010101101101100;
   assign mem[11030] = 32'b11111011011011101100111111100000;
   assign mem[11031] = 32'b00000001011001110000011110010100;
   assign mem[11032] = 32'b00000000010010000110000010001000;
   assign mem[11033] = 32'b11111011000110001010000010000000;
   assign mem[11034] = 32'b11111111110001010110011101111011;
   assign mem[11035] = 32'b11111100101001000101111001001100;
   assign mem[11036] = 32'b11110101000100100000101010110000;
   assign mem[11037] = 32'b11111111110100011001001000111010;
   assign mem[11038] = 32'b00000100001001001111100100001000;
   assign mem[11039] = 32'b00000000110010101100111010011100;
   assign mem[11040] = 32'b11111111011110000110100110100010;
   assign mem[11041] = 32'b11111100100001010101001110000000;
   assign mem[11042] = 32'b00000010101011001110001101011100;
   assign mem[11043] = 32'b00000100011111010011100000100000;
   assign mem[11044] = 32'b11111111100000001110110110011111;
   assign mem[11045] = 32'b00000011100001110110001110011100;
   assign mem[11046] = 32'b00000000110111100011001111000000;
   assign mem[11047] = 32'b11111001001001101101101101011000;
   assign mem[11048] = 32'b00000010000011111011111110001000;
   assign mem[11049] = 32'b00000011010111001000010011101000;
   assign mem[11050] = 32'b11110110110011111001001011110000;
   assign mem[11051] = 32'b00000001010010110111100011110100;
   assign mem[11052] = 32'b11111100011111011100001000101100;
   assign mem[11053] = 32'b11111011111101101110000100110000;
   assign mem[11054] = 32'b00000001101100011100100000000010;
   assign mem[11055] = 32'b11111101100000011111101001001100;
   assign mem[11056] = 32'b00000010010110001100000000010000;
   assign mem[11057] = 32'b00000011110110101110101001000100;
   assign mem[11058] = 32'b11111100011111100100010111000000;
   assign mem[11059] = 32'b00000101101101010010000110111000;
   assign mem[11060] = 32'b11111011011011110010111111011000;
   assign mem[11061] = 32'b00000101110110101101111011010000;
   assign mem[11062] = 32'b11111010111001010111011110011000;
   assign mem[11063] = 32'b00000100001101010101101011111000;
   assign mem[11064] = 32'b00000000100010111100011010010011;
   assign mem[11065] = 32'b00000010010001111000111110010100;
   assign mem[11066] = 32'b00000000110111000100111001000111;
   assign mem[11067] = 32'b11111000000100001100000010111000;
   assign mem[11068] = 32'b11111100000110001001111010011100;
   assign mem[11069] = 32'b00000001001011101111000110110110;
   assign mem[11070] = 32'b00000011011001110100000101101000;
   assign mem[11071] = 32'b11101100110110110011101011100000;
   assign mem[11072] = 32'b00000011010101000011010101011100;
   assign mem[11073] = 32'b00000011100000110010001001101000;
   assign mem[11074] = 32'b00000010001100111110101101010000;
   assign mem[11075] = 32'b11111111000001000000000001010000;
   assign mem[11076] = 32'b00000000000111110001111100101111;
   assign mem[11077] = 32'b11111010001000001010000111110000;
   assign mem[11078] = 32'b11111110000110001010000000101110;
   assign mem[11079] = 32'b00001000000011100011110001100000;
   assign mem[11080] = 32'b11110110001011001000010001000000;
   assign mem[11081] = 32'b00000100101110000101111100011000;
   assign mem[11082] = 32'b11111011110100011000010100001000;
   assign mem[11083] = 32'b11111100001111010110110011101100;
   assign mem[11084] = 32'b11111111011000000001100101110110;
   assign mem[11085] = 32'b11111010110011010010010000111000;
   assign mem[11086] = 32'b11111011100101111011010000001000;
   assign mem[11087] = 32'b00000010010100000001001100111100;
   assign mem[11088] = 32'b00000000001101010000001111010010;
   assign mem[11089] = 32'b00000011110111011100001000101000;
   assign mem[11090] = 32'b00000000111010111101000010011110;
   assign mem[11091] = 32'b11111000110011110010001000111000;
   assign mem[11092] = 32'b11111101110010011000000011111100;
   assign mem[11093] = 32'b11111111100100100011001110010010;
   assign mem[11094] = 32'b11111100010001010000100101010000;
   assign mem[11095] = 32'b11111101110111111001100111100100;
   assign mem[11096] = 32'b11111011110000100110001101111000;
   assign mem[11097] = 32'b00000001110010111011101001000000;
   assign mem[11098] = 32'b11111110100010011001000110011110;
   assign mem[11099] = 32'b00000001001110010110011001100000;
   assign mem[11100] = 32'b00000011001011111001000100110100;
   assign mem[11101] = 32'b11111111100011010000011001010101;
   assign mem[11102] = 32'b00000011001000010011110000100100;
   assign mem[11103] = 32'b11111000000110011010011101111000;
   assign mem[11104] = 32'b11111111011011110011000101000011;
   assign mem[11105] = 32'b11111011000001101110100111111000;
   assign mem[11106] = 32'b11111001100001000010100000010000;
   assign mem[11107] = 32'b11111111010001001011100111100110;
   assign mem[11108] = 32'b00000100101111100110101000110000;
   assign mem[11109] = 32'b00000010000111000001011010111000;
   assign mem[11110] = 32'b00000111100111000111110000000000;
   assign mem[11111] = 32'b00000100110000010110111111110000;
   assign mem[11112] = 32'b11111010001110011110011001111000;
   assign mem[11113] = 32'b00000100111110010001010000010000;
   assign mem[11114] = 32'b11111011010000100100100110010000;
   assign mem[11115] = 32'b11111111111001011011110110001000;
   assign mem[11116] = 32'b00000011000111110101000110101100;
   assign mem[11117] = 32'b11111001011001001010011100010000;
   assign mem[11118] = 32'b00000010110100100100001110111100;
   assign mem[11119] = 32'b11111001111001101001100111100000;
   assign mem[11120] = 32'b00000111111100010101100100010000;
   assign mem[11121] = 32'b00001001100010100110001010000000;
   assign mem[11122] = 32'b11110101011010101011010011000000;
   assign mem[11123] = 32'b00000101000001111100010001101000;
   assign mem[11124] = 32'b11110111000111011101110111100000;
   assign mem[11125] = 32'b00000110011100111011101111100000;
   assign mem[11126] = 32'b00000111010010011001100101110000;
   assign mem[11127] = 32'b11110001001000011001100000000000;
   assign mem[11128] = 32'b00000011101011111100001011001100;
   assign mem[11129] = 32'b11111010010100001100100001011000;
   assign mem[11130] = 32'b00000100111011100101100110000000;
   assign mem[11131] = 32'b00001100110110110001001010100000;
   assign mem[11132] = 32'b00000011000101100110010110101000;
   assign mem[11133] = 32'b11110101110111000110010001110000;
   assign mem[11134] = 32'b11110111100001111010101011010000;
   assign mem[11135] = 32'b11111011100001011010010010011000;
   assign mem[11136] = 32'b11111101100100010100100110100000;
   assign mem[11137] = 32'b00001011101100111100010001110000;
   assign mem[11138] = 32'b11111111110000101101000000001111;
   assign mem[11139] = 32'b11101101100010011001110100100000;
   assign mem[11140] = 32'b00000110110100000001001100111000;
   assign mem[11141] = 32'b11111111001110100011101001011000;
   assign mem[11142] = 32'b00000001000001111001010110101000;
   assign mem[11143] = 32'b11110001101010101011010111100000;
   assign mem[11144] = 32'b00000000010101010000100001001011;
   assign mem[11145] = 32'b00000000110111101010111110001101;
   assign mem[11146] = 32'b00000011110001011100001011110000;
   assign mem[11147] = 32'b11111011111011000101110111101000;
   assign mem[11148] = 32'b00000010110000100111111011010000;
   assign mem[11149] = 32'b11111010001001010011100011010000;
   assign mem[11150] = 32'b00000001110011000100001100010000;
   assign mem[11151] = 32'b00000100000011010001100010110000;
   assign mem[11152] = 32'b00000101001101011011011100110000;
   assign mem[11153] = 32'b11111010110011010110011001110000;
   assign mem[11154] = 32'b11111100000100011110000111110100;
   assign mem[11155] = 32'b11111101100111101010101010001000;
   assign mem[11156] = 32'b11111110101000011001100100010110;
   assign mem[11157] = 32'b00001001101111010010000100000000;
   assign mem[11158] = 32'b11111001110101011111111101011000;
   assign mem[11159] = 32'b11111001001011001000101101010000;
   assign mem[11160] = 32'b00000010001101011100101011010100;
   assign mem[11161] = 32'b11111001000001011111111111100000;
   assign mem[11162] = 32'b00000010110011100110110110101100;
   assign mem[11163] = 32'b11111011110100110001110010100000;
   assign mem[11164] = 32'b00000101111000111110101101001000;
   assign mem[11165] = 32'b11111111001101110010010101010010;
   assign mem[11166] = 32'b11111101101011000000001110100100;
   assign mem[11167] = 32'b11111010000010000111001101000000;
   assign mem[11168] = 32'b00000000010101001000001001101110;
   assign mem[11169] = 32'b00001001000100111010100101000000;
   assign mem[11170] = 32'b00000011111010110100100100111100;
   assign mem[11171] = 32'b00001011101100100000100000100000;
   assign mem[11172] = 32'b00000000010010101010111110100101;
   assign mem[11173] = 32'b00000010000000101011101011010100;
   assign mem[11174] = 32'b00000101000010111100110110101000;
   assign mem[11175] = 32'b00000000000110100001110101110010;
   assign mem[11176] = 32'b11111110000110010101111011100110;
   assign mem[11177] = 32'b00001000110010111000101011000000;
   assign mem[11178] = 32'b11110010111000111011100110100000;
   assign mem[11179] = 32'b11111100011011110101011011000000;
   assign mem[11180] = 32'b00000101000000100001000011000000;
   assign mem[11181] = 32'b00000011010000001110010110011000;
   assign mem[11182] = 32'b11111111010011011010010000110111;
   assign mem[11183] = 32'b11110111100111110100011110000000;
   assign mem[11184] = 32'b11111111000110101100101111110101;
   assign mem[11185] = 32'b11111111101110010110111101001000;
   assign mem[11186] = 32'b00000101110111100001011001000000;
   assign mem[11187] = 32'b11111110000111101110011101001000;
   assign mem[11188] = 32'b00000000110111001011110011011010;
   assign mem[11189] = 32'b00000000001011101010000101001111;
   assign mem[11190] = 32'b11111100110111111000100000011100;
   assign mem[11191] = 32'b11111001111000001110101010101000;
   assign mem[11192] = 32'b11111111010101001011101111000100;
   assign mem[11193] = 32'b00000010110110000011010010001100;
   assign mem[11194] = 32'b00000100100101101101100100111000;
   assign mem[11195] = 32'b00000001011001011100101000000100;
   assign mem[11196] = 32'b00000001010011001110000111101010;
   assign mem[11197] = 32'b11111111001001010101100101010110;
   assign mem[11198] = 32'b11111011000101000111111111011000;
   assign mem[11199] = 32'b00000100001111110001000100110000;
   assign mem[11200] = 32'b11111001010111100110000100011000;
   assign mem[11201] = 32'b11111110000001101101111000111010;
   assign mem[11202] = 32'b00000100000001000011011000011000;
   assign mem[11203] = 32'b11111111101000110010110100010001;
   assign mem[11204] = 32'b11111001100100011001010101100000;
   assign mem[11205] = 32'b11111110001010100100010101010100;
   assign mem[11206] = 32'b00000010001001011110001111111100;
   assign mem[11207] = 32'b00000010100111011100100001001000;
   assign mem[11208] = 32'b00000011011000100111101111001100;
   assign mem[11209] = 32'b11111111001011101010001101011101;
   assign mem[11210] = 32'b11111111100111101010010000011010;
   assign mem[11211] = 32'b00000101100000111011011010101000;
   assign mem[11212] = 32'b00000101001110010110010010111000;
   assign mem[11213] = 32'b11111011000000100100000101011000;
   assign mem[11214] = 32'b00000010011010000011011011011100;
   assign mem[11215] = 32'b00000100100111111101111101111000;
   assign mem[11216] = 32'b11111111110010111011000001011011;
   assign mem[11217] = 32'b00000010001100010010011100110000;
   assign mem[11218] = 32'b11111001010100111101111110101000;
   assign mem[11219] = 32'b11111111010101101011100000110001;
   assign mem[11220] = 32'b11111010000010110100110011010000;
   assign mem[11221] = 32'b11111101000000011010110001110100;
   assign mem[11222] = 32'b00000000101110000111000000110100;
   assign mem[11223] = 32'b00000000110001001110100001110101;
   assign mem[11224] = 32'b00000110011011100101101101110000;
   assign mem[11225] = 32'b00000000000111011101111000110100;
   assign mem[11226] = 32'b11111111100100100001100110000101;
   assign mem[11227] = 32'b11111011110101010111100111000000;
   assign mem[11228] = 32'b11111110001110101011000000101010;
   assign mem[11229] = 32'b00000000001000111010100111101001;
   assign mem[11230] = 32'b00001010100001111001110011110000;
   assign mem[11231] = 32'b00011000001110101100011010100000;
   assign mem[11232] = 32'b00000010000110011110111101001000;
   assign mem[11233] = 32'b11111100010010011100110000010100;
   assign mem[11234] = 32'b11110001001110110000001110010000;
   assign mem[11235] = 32'b11111110101110010011101101101110;
   assign mem[11236] = 32'b11111101111001111111111100011100;
   assign mem[11237] = 32'b00001110011010011000010010000000;
   assign mem[11238] = 32'b11111000110010011011100010010000;
   assign mem[11239] = 32'b11101111111101111010101111100000;
   assign mem[11240] = 32'b00000100110110111010001110000000;
   assign mem[11241] = 32'b11111010100100110100101110011000;
   assign mem[11242] = 32'b11111011100001011101101011001000;
   assign mem[11243] = 32'b00001000010000001001100001100000;
   assign mem[11244] = 32'b11111111011110011100001001010101;
   assign mem[11245] = 32'b00000010110100010110001001010000;
   assign mem[11246] = 32'b11111010010010111010011101101000;
   assign mem[11247] = 32'b11111000110010001011010000000000;
   assign mem[11248] = 32'b11111101110011001000110000000100;
   assign mem[11249] = 32'b00000010101000111000000110011100;
   assign mem[11250] = 32'b00000011101001000111111110011000;
   assign mem[11251] = 32'b11110010100110000110100001100000;
   assign mem[11252] = 32'b00000010001010001011100110110000;
   assign mem[11253] = 32'b11111101000111111011000001110100;
   assign mem[11254] = 32'b11111111101011000011111010011110;
   assign mem[11255] = 32'b00000110111011101100100101110000;
   assign mem[11256] = 32'b00000011011000011101010011100000;
   assign mem[11257] = 32'b11110111101001011010101100010000;
   assign mem[11258] = 32'b11111001011111011111101011001000;
   assign mem[11259] = 32'b00000001011111010110001100100000;
   assign mem[11260] = 32'b11111110000001001000101111000100;
   assign mem[11261] = 32'b11110111101011011000001001110000;
   assign mem[11262] = 32'b00000010001010001101100000100000;
   assign mem[11263] = 32'b11111100111011010101011010100100;
   assign mem[11264] = 32'b00000101101100011000000011010000;
   assign mem[11265] = 32'b00000010001111001100011010000100;
   assign mem[11266] = 32'b11111111101000111000101001000010;
   assign mem[11267] = 32'b11110001110101101000000000010000;
   assign mem[11268] = 32'b11111110011101011101111011100110;
   assign mem[11269] = 32'b00000110110000000110011011011000;
   assign mem[11270] = 32'b11111010100010101110100110011000;
   assign mem[11271] = 32'b11110100100101110101100001000000;
   assign mem[11272] = 32'b11110101111011100010011111110000;
   assign mem[11273] = 32'b00000111110101100011011000100000;
   assign mem[11274] = 32'b00000100011001111101000100101000;
   assign mem[11275] = 32'b00000001111100111111100110110110;
   assign mem[11276] = 32'b11110101000110000011010010000000;
   assign mem[11277] = 32'b00000001101110110010011111000010;
   assign mem[11278] = 32'b11111010010101010110111001100000;
   assign mem[11279] = 32'b00001000100000010111111000010000;
   assign mem[11280] = 32'b11110100011110110101101011110000;
   assign mem[11281] = 32'b00000111101000110111100110100000;
   assign mem[11282] = 32'b00000100000001001101001100010000;
   assign mem[11283] = 32'b00000110001100111000011001000000;
   assign mem[11284] = 32'b00000000011000101101001111010101;
   assign mem[11285] = 32'b00000001000111100101000110111010;
   assign mem[11286] = 32'b11111100010011101110100000011000;
   assign mem[11287] = 32'b11111000011001101000101110011000;
   assign mem[11288] = 32'b00000000100111001110100000101111;
   assign mem[11289] = 32'b11111101110001010101010010000100;
   assign mem[11290] = 32'b11101100101001100101010010100000;
   assign mem[11291] = 32'b00000110101000101100001101000000;
   assign mem[11292] = 32'b00000001010100000110101111001000;
   assign mem[11293] = 32'b00000011101011100100001011001100;
   assign mem[11294] = 32'b00000010100100001010111010110000;
   assign mem[11295] = 32'b00000011100111100111100011100100;
   assign mem[11296] = 32'b11111010101111110000010111111000;
   assign mem[11297] = 32'b11111011010101010100010101001000;
   assign mem[11298] = 32'b11111110010111001011100101001000;
   assign mem[11299] = 32'b00000101001100000111000110000000;
   assign mem[11300] = 32'b11111000000000111100110100111000;
   assign mem[11301] = 32'b11110100111110000000110100000000;
   assign mem[11302] = 32'b11111001101101100001001101001000;
   assign mem[11303] = 32'b00001011001110111111010000010000;
   assign mem[11304] = 32'b00000100000101001000000110110000;
   assign mem[11305] = 32'b00000001110100011100100110011110;
   assign mem[11306] = 32'b11111011000110110000111110000000;
   assign mem[11307] = 32'b11111000111011000110110000100000;
   assign mem[11308] = 32'b11110110110010010110111000000000;
   assign mem[11309] = 32'b00000110100010011101111001111000;
   assign mem[11310] = 32'b00001000110111000100011010100000;
   assign mem[11311] = 32'b00000010001011000111010111110000;
   assign mem[11312] = 32'b00000001100100001110111011000010;
   assign mem[11313] = 32'b00000011100001101010101000110000;
   assign mem[11314] = 32'b11110111111101111110001000110000;
   assign mem[11315] = 32'b00000000111100000010001001011001;
   assign mem[11316] = 32'b00000110000110000001011011111000;
   assign mem[11317] = 32'b11111011010010110001011000001000;
   assign mem[11318] = 32'b00000111100001110001100000001000;
   assign mem[11319] = 32'b11101111111011110101111101000000;
   assign mem[11320] = 32'b11111100100111010010110010001000;
   assign mem[11321] = 32'b11111100011001001101001101011000;
   assign mem[11322] = 32'b00000011101011000111110111110100;
   assign mem[11323] = 32'b00000011101110110010001111001000;
   assign mem[11324] = 32'b00000111010101001010111100011000;
   assign mem[11325] = 32'b11111111101001110010100111100110;
   assign mem[11326] = 32'b00001001110101010111110010110000;
   assign mem[11327] = 32'b11111011011111110101100011101000;
   assign mem[11328] = 32'b11111000101110110010011011100000;
   assign mem[11329] = 32'b11111110001010100110110111010100;
   assign mem[11330] = 32'b11110100010100010111011010110000;
   assign mem[11331] = 32'b00000011001000000101010010110000;
   assign mem[11332] = 32'b11111110110001001100111010000010;
   assign mem[11333] = 32'b11111101110110101010101110010000;
   assign mem[11334] = 32'b00000011110011010001000011100000;
   assign mem[11335] = 32'b00000101011101000011011011101000;
   assign mem[11336] = 32'b00000000111011101101101110010100;
   assign mem[11337] = 32'b11111010111100111100001010101000;
   assign mem[11338] = 32'b00000110010010100101110010011000;
   assign mem[11339] = 32'b11111010010010011011110010011000;
   assign mem[11340] = 32'b11101010010100111101101000100000;
   assign mem[11341] = 32'b00001100100100000110101011110000;
   assign mem[11342] = 32'b11111100010000110100101000000000;
   assign mem[11343] = 32'b11111011101011111101101100010000;
   assign mem[11344] = 32'b00001000011100010110100000010000;
   assign mem[11345] = 32'b11111111010000110000000100111110;
   assign mem[11346] = 32'b11110111110101111011010101110000;
   assign mem[11347] = 32'b00000001001101000010011010111000;
   assign mem[11348] = 32'b11111101100101100110111111000100;
   assign mem[11349] = 32'b00000011101111101001011001101100;
   assign mem[11350] = 32'b11111100110111111001010001011000;
   assign mem[11351] = 32'b00000001100001100101011001100110;
   assign mem[11352] = 32'b11111111101110001000100011110111;
   assign mem[11353] = 32'b11111111101100011000001010011110;
   assign mem[11354] = 32'b11111101101111011011011010011100;
   assign mem[11355] = 32'b11111111101101111111011100010110;
   assign mem[11356] = 32'b00000001100110100110010000100110;
   assign mem[11357] = 32'b00000000010011100111001010011011;
   assign mem[11358] = 32'b11111011111000111011010010010000;
   assign mem[11359] = 32'b00000010011001011000101010101000;
   assign mem[11360] = 32'b11110011010010110110100001110000;
   assign mem[11361] = 32'b00000100110110101000101001110000;
   assign mem[11362] = 32'b00000101010100100011001000100000;
   assign mem[11363] = 32'b11111011101100010101001110000000;
   assign mem[11364] = 32'b11111010011011100100011000111000;
   assign mem[11365] = 32'b11111011000001100000111011110000;
   assign mem[11366] = 32'b00000000001100000011010011101001;
   assign mem[11367] = 32'b00000101011110010111010000001000;
   assign mem[11368] = 32'b00000011111101101111111011011100;
   assign mem[11369] = 32'b11110100011001010100111010000000;
   assign mem[11370] = 32'b11111100010100101010010001000100;
   assign mem[11371] = 32'b00000010000111001001000010000100;
   assign mem[11372] = 32'b00000010011110110011110001010100;
   assign mem[11373] = 32'b11111110101000001101010011101100;
   assign mem[11374] = 32'b00000001101010010011000000000000;
   assign mem[11375] = 32'b11111101011111110101101101111100;
   assign mem[11376] = 32'b00000000100111001000011110110111;
   assign mem[11377] = 32'b11111111000000000110111111111101;
   assign mem[11378] = 32'b11111101010000101110001100011100;
   assign mem[11379] = 32'b11111101111110011111101001001000;
   assign mem[11380] = 32'b00001000011011011110100110000000;
   assign mem[11381] = 32'b11111000000011010100010110111000;
   assign mem[11382] = 32'b00000010100110010101000000100000;
   assign mem[11383] = 32'b11111101000011010111100100110100;
   assign mem[11384] = 32'b00000000110000101010001101011110;
   assign mem[11385] = 32'b11111100011111110111000111010100;
   assign mem[11386] = 32'b00000000010100110000011111110100;
   assign mem[11387] = 32'b11111111001101101011000110011010;
   assign mem[11388] = 32'b00000001001000001010001010001010;
   assign mem[11389] = 32'b00000011001100001011111100101000;
   assign mem[11390] = 32'b11110000001011011110111110110000;
   assign mem[11391] = 32'b00001011111100101111110111010000;
   assign mem[11392] = 32'b11110100100100001111111011110000;
   assign mem[11393] = 32'b00000101001001110111101101110000;
   assign mem[11394] = 32'b00000010011010000000000100000000;
   assign mem[11395] = 32'b00000011010011010010010110010000;
   assign mem[11396] = 32'b11111010111101110110000000001000;
   assign mem[11397] = 32'b00000011011110100010110110100000;
   assign mem[11398] = 32'b11110001011000110000000100100000;
   assign mem[11399] = 32'b00000100101011101000001110001000;
   assign mem[11400] = 32'b11111101010001001011101001101100;
   assign mem[11401] = 32'b11110110010000101011000001010000;
   assign mem[11402] = 32'b11111010111010001001110011010000;
   assign mem[11403] = 32'b00000000111001111000100011110110;
   assign mem[11404] = 32'b00000010011100100101101000101100;
   assign mem[11405] = 32'b11111100111011101110001000110100;
   assign mem[11406] = 32'b11111110001100101000000110001010;
   assign mem[11407] = 32'b00000000101111101011010111010110;
   assign mem[11408] = 32'b11111101011000111011010110111100;
   assign mem[11409] = 32'b00000100100011111100010111110000;
   assign mem[11410] = 32'b11111110010100101000010001101000;
   assign mem[11411] = 32'b11110100110001001001100110100000;
   assign mem[11412] = 32'b11111110010100011011111111101110;
   assign mem[11413] = 32'b00000100011011100110101001010000;
   assign mem[11414] = 32'b00000100111000100011001100000000;
   assign mem[11415] = 32'b00000000011010111001011010110000;
   assign mem[11416] = 32'b11111111000011101110000000011101;
   assign mem[11417] = 32'b11111111110111001110000101101010;
   assign mem[11418] = 32'b11111000101011000100100110111000;
   assign mem[11419] = 32'b11111110110010001010101101001110;
   assign mem[11420] = 32'b00000000100100001100001011001100;
   assign mem[11421] = 32'b00000001010011101011111000010010;
   assign mem[11422] = 32'b00000010110111111110101010000100;
   assign mem[11423] = 32'b00000111111001101110101001110000;
   assign mem[11424] = 32'b11111011110100101001110111001000;
   assign mem[11425] = 32'b11111011011100000100011111110000;
   assign mem[11426] = 32'b00000000000010100000000110011111;
   assign mem[11427] = 32'b11111101111010011101100010100000;
   assign mem[11428] = 32'b11111111100101010000000101001001;
   assign mem[11429] = 32'b11111100011110000100111011111100;
   assign mem[11430] = 32'b00001111100010011111110111010000;
   assign mem[11431] = 32'b00000001110011010111101001110100;
   assign mem[11432] = 32'b11111111010001101011101011001001;
   assign mem[11433] = 32'b11101110111110010101011111000000;
   assign mem[11434] = 32'b11111001000101101111001000100000;
   assign mem[11435] = 32'b00000000001111001101010010110100;
   assign mem[11436] = 32'b11111101010011111010110011001000;
   assign mem[11437] = 32'b00000000101001010110111010010111;
   assign mem[11438] = 32'b00000011010010000100010101000000;
   assign mem[11439] = 32'b11111001010011001101010011111000;
   assign mem[11440] = 32'b00000000110110111101001100011010;
   assign mem[11441] = 32'b00001100000101101000001101100000;
   assign mem[11442] = 32'b11111011110010011101011001001000;
   assign mem[11443] = 32'b00000110001001110010010100010000;
   assign mem[11444] = 32'b00000000111111011111110110101101;
   assign mem[11445] = 32'b00000001001011100001101111011000;
   assign mem[11446] = 32'b00000100101101010100100110001000;
   assign mem[11447] = 32'b11111011010110001011000010000000;
   assign mem[11448] = 32'b11111101011010110110111010100100;
   assign mem[11449] = 32'b11110100001100101110101011000000;
   assign mem[11450] = 32'b11110001001001000001011010110000;
   assign mem[11451] = 32'b11111010010110111010011110010000;
   assign mem[11452] = 32'b11111110110011110010011100011110;
   assign mem[11453] = 32'b00000000001101010111011111000101;
   assign mem[11454] = 32'b00001000101001111010111010000000;
   assign mem[11455] = 32'b00000011100000001100110110110000;
   assign mem[11456] = 32'b11111000011111001001111000001000;
   assign mem[11457] = 32'b11111010110011111000100000001000;
   assign mem[11458] = 32'b11111111100100110101001110101101;
   assign mem[11459] = 32'b00000011001100111100111011110100;
   assign mem[11460] = 32'b00000101100101100111100110110000;
   assign mem[11461] = 32'b00000010101011000111011011101000;
   assign mem[11462] = 32'b00000010010011000110100011010100;
   assign mem[11463] = 32'b00000101101000001101011110001000;
   assign mem[11464] = 32'b11111101000011010111110000100100;
   assign mem[11465] = 32'b00000001000110001000010100100110;
   assign mem[11466] = 32'b11111010110000011101110101110000;
   assign mem[11467] = 32'b11111010111011100010111000101000;
   assign mem[11468] = 32'b11110000010000001111001110110000;
   assign mem[11469] = 32'b11111110101100101011101110110000;
   assign mem[11470] = 32'b11111101000011111110000000100100;
   assign mem[11471] = 32'b00000100101111011010101100011000;
   assign mem[11472] = 32'b00000001010010011000010111111100;
   assign mem[11473] = 32'b00000011001000011110011100000100;
   assign mem[11474] = 32'b11111011010110101011100000000000;
   assign mem[11475] = 32'b00000010101011101001000110000100;
   assign mem[11476] = 32'b00001000010010011101011011010000;
   assign mem[11477] = 32'b11111010011101101101011010101000;
   assign mem[11478] = 32'b00001001000111101011111000100000;
   assign mem[11479] = 32'b11110110010111010110010100110000;
   assign mem[11480] = 32'b00000011010101001001111001101000;
   assign mem[11481] = 32'b11111100000101110101010011001000;
   assign mem[11482] = 32'b00000101100101111000110000111000;
   assign mem[11483] = 32'b11111111110100101001010110001110;
   assign mem[11484] = 32'b11111011000001010111010011111000;
   assign mem[11485] = 32'b00000011110011000010001111010100;
   assign mem[11486] = 32'b11110110000111000100000100010000;
   assign mem[11487] = 32'b00000101010011101001001110001000;
   assign mem[11488] = 32'b11111000110100000101001110011000;
   assign mem[11489] = 32'b00000001001111111110110000010100;
   assign mem[11490] = 32'b11111111011101101011010100110010;
   assign mem[11491] = 32'b00000010000101011001111011100000;
   assign mem[11492] = 32'b00000101100000010100010011101000;
   assign mem[11493] = 32'b11111110001011010111110010000100;
   assign mem[11494] = 32'b11111100100001111101000101111100;
   assign mem[11495] = 32'b00000000111001011000101111100000;
   assign mem[11496] = 32'b00000011001111100100111100011100;
   assign mem[11497] = 32'b00000000100010001110000010101000;
   assign mem[11498] = 32'b11111111100110001001101100100100;
   assign mem[11499] = 32'b00000011111010110001011011010000;
   assign mem[11500] = 32'b11110101111011011110001001010000;
   assign mem[11501] = 32'b00000111101011101000110100111000;
   assign mem[11502] = 32'b11111001110011110010000011011000;
   assign mem[11503] = 32'b00000001010101110010010110111010;
   assign mem[11504] = 32'b11110111110101000011000010100000;
   assign mem[11505] = 32'b00000001111111010010100010001010;
   assign mem[11506] = 32'b11111111110111111110111111000001;
   assign mem[11507] = 32'b00000010011111111001101111100000;
   assign mem[11508] = 32'b11111001101111000001111100010000;
   assign mem[11509] = 32'b11111111101010001100111000011001;
   assign mem[11510] = 32'b11111100100000010110000100011100;
   assign mem[11511] = 32'b00000111010011101011111010101000;
   assign mem[11512] = 32'b00000101000111100101110100001000;
   assign mem[11513] = 32'b11111101110000111001001001001000;
   assign mem[11514] = 32'b11111110101101100101110110101000;
   assign mem[11515] = 32'b11111111010011111111000000010011;
   assign mem[11516] = 32'b00000100001101101000111100011000;
   assign mem[11517] = 32'b11111111100000110010111110000010;
   assign mem[11518] = 32'b11111011101101000001001101001000;
   assign mem[11519] = 32'b11111110010111011010100101101000;
   assign mem[11520] = 32'b00000010001010000011001101011100;
   assign mem[11521] = 32'b11110110011110001101010011100000;
   assign mem[11522] = 32'b00000010010000101000000101110100;
   assign mem[11523] = 32'b11111111100101000001001011100010;
   assign mem[11524] = 32'b11111101010000101000110011111000;
   assign mem[11525] = 32'b00000000010000001101000111001111;
   assign mem[11526] = 32'b00000000101001011011011011011111;
   assign mem[11527] = 32'b00000001101100000001110001110110;
   assign mem[11528] = 32'b00000111010011001101011010110000;
   assign mem[11529] = 32'b11111000101000011000101100111000;
   assign mem[11530] = 32'b11111100100111111010010111011100;
   assign mem[11531] = 32'b00000001111001010101100000111100;
   assign mem[11532] = 32'b11110100101100101110101100110000;
   assign mem[11533] = 32'b00000011111101100110010110001000;
   assign mem[11534] = 32'b11101000010010011010000101000000;
   assign mem[11535] = 32'b00000111111001111000000011111000;
   assign mem[11536] = 32'b00001100111001100101001011000000;
   assign mem[11537] = 32'b11110000100111111100011000100000;
   assign mem[11538] = 32'b00000010000000010001000000111100;
   assign mem[11539] = 32'b11111001011001111001011100110000;
   assign mem[11540] = 32'b11110111100011010101001000110000;
   assign mem[11541] = 32'b11111110010011110001110010010100;
   assign mem[11542] = 32'b00000101011110000110000011011000;
   assign mem[11543] = 32'b00000110110100110000000101011000;
   assign mem[11544] = 32'b11111001011000100000100100111000;
   assign mem[11545] = 32'b00000111011001010010100100011000;
   assign mem[11546] = 32'b00000001001010110010010110101110;
   assign mem[11547] = 32'b11110101000001000110011111000000;
   assign mem[11548] = 32'b00000010001100000101111110111000;
   assign mem[11549] = 32'b11110101000111101110011111100000;
   assign mem[11550] = 32'b11111110000001010111111011010100;
   assign mem[11551] = 32'b11110011000101011100000001000000;
   assign mem[11552] = 32'b00000000100111001011111010001110;
   assign mem[11553] = 32'b00000011111101111101110111110100;
   assign mem[11554] = 32'b11111101101011000110100101111000;
   assign mem[11555] = 32'b11111111010000100010000001010000;
   assign mem[11556] = 32'b11111110110111001111010111010000;
   assign mem[11557] = 32'b11111100000101000101000101011000;
   assign mem[11558] = 32'b11111101011001110111011011001100;
   assign mem[11559] = 32'b11111110001101001011111000011000;
   assign mem[11560] = 32'b00000000101101010001000001101010;
   assign mem[11561] = 32'b00001000111011011101001001010000;
   assign mem[11562] = 32'b11111101010111001101100110111100;
   assign mem[11563] = 32'b00000000010001110100111000010001;
   assign mem[11564] = 32'b11111101101011111011010011111000;
   assign mem[11565] = 32'b11110111101110100011000100110000;
   assign mem[11566] = 32'b11110111001010011000101100110000;
   assign mem[11567] = 32'b00000010110100001000010011001100;
   assign mem[11568] = 32'b00000101111110111001000011001000;
   assign mem[11569] = 32'b11111110100101011010110011111010;
   assign mem[11570] = 32'b11111111101001010011111111000100;
   assign mem[11571] = 32'b00000001111110110000101000100100;
   assign mem[11572] = 32'b00000010101001001100100111010100;
   assign mem[11573] = 32'b11111101010110001001100011010000;
   assign mem[11574] = 32'b11111011111010011110011001100000;
   assign mem[11575] = 32'b00000010000011011001000010011000;
   assign mem[11576] = 32'b00000001010000000100101010100110;
   assign mem[11577] = 32'b00000100010001011011110010111000;
   assign mem[11578] = 32'b11111000011000011000000111001000;
   assign mem[11579] = 32'b11111111011110000100100011011000;
   assign mem[11580] = 32'b11111010111010111011100011011000;
   assign mem[11581] = 32'b00000100111101111000111010110000;
   assign mem[11582] = 32'b11111110011101010101100000011100;
   assign mem[11583] = 32'b00000001111011100110011110001010;
   assign mem[11584] = 32'b11111011111110101000010101011000;
   assign mem[11585] = 32'b00000001011010001101001101011110;
   assign mem[11586] = 32'b11111010111101011000000011101000;
   assign mem[11587] = 32'b11111111100010000100100111000101;
   assign mem[11588] = 32'b11111110101010011011111111001000;
   assign mem[11589] = 32'b00000001100001011000110011000010;
   assign mem[11590] = 32'b00000101111100011010001111010000;
   assign mem[11591] = 32'b11111010100010010100101001101000;
   assign mem[11592] = 32'b00000001001101011110011000000000;
   assign mem[11593] = 32'b00000011010001010001101010010000;
   assign mem[11594] = 32'b11111011011101100010000101110000;
   assign mem[11595] = 32'b11111100010001110101010000011000;
   assign mem[11596] = 32'b00000000110010110011000011111101;
   assign mem[11597] = 32'b00000000111101001011001010010001;
   assign mem[11598] = 32'b00000100101000011111111110110000;
   assign mem[11599] = 32'b00000000101111111100100001001011;
   assign mem[11600] = 32'b00010000101000000111011011100000;
   assign mem[11601] = 32'b11110010001110010101000111110000;
   assign mem[11602] = 32'b00000010011110010100101010011000;
   assign mem[11603] = 32'b11111100010011101000100000101000;
   assign mem[11604] = 32'b11110100011011000001000100010000;
   assign mem[11605] = 32'b00000010011001100111100111101000;
   assign mem[11606] = 32'b00000010010101010011101111101100;
   assign mem[11607] = 32'b00000101110010000001011001110000;
   assign mem[11608] = 32'b11111001011110101010000111101000;
   assign mem[11609] = 32'b11110000000101110011100101010000;
   assign mem[11610] = 32'b00000001000111100011010110000010;
   assign mem[11611] = 32'b00010110100101011000001000100000;
   assign mem[11612] = 32'b11110101011100000110100011100000;
   assign mem[11613] = 32'b00000001000110011010010100010010;
   assign mem[11614] = 32'b11111111101010110111101100101001;
   assign mem[11615] = 32'b00001000110111010101011000110000;
   assign mem[11616] = 32'b11110110011010010011011000000000;
   assign mem[11617] = 32'b00001000001010110111101011100000;
   assign mem[11618] = 32'b11110101011000011011111011010000;
   assign mem[11619] = 32'b11111101010100111001101101000100;
   assign mem[11620] = 32'b00000011001001111100000010011000;
   assign mem[11621] = 32'b11111010100000000110110100000000;
   assign mem[11622] = 32'b00000001000101100110010100100110;
   assign mem[11623] = 32'b11111000010100011000010110101000;
   assign mem[11624] = 32'b00000001100010010111111001010000;
   assign mem[11625] = 32'b11111110001010110011100010001100;
   assign mem[11626] = 32'b00000000100011001110000101111101;
   assign mem[11627] = 32'b00000010000011110111000011101100;
   assign mem[11628] = 32'b00001001001011101111001111110000;
   assign mem[11629] = 32'b00000100110010110011010110010000;
   assign mem[11630] = 32'b00000001010110000001000110110010;
   assign mem[11631] = 32'b11111100001001101100000111101100;
   assign mem[11632] = 32'b11111110001110111001000110010000;
   assign mem[11633] = 32'b00000101101010010010011110101000;
   assign mem[11634] = 32'b11111101100110110000011010010100;
   assign mem[11635] = 32'b00000110001000100000101100110000;
   assign mem[11636] = 32'b00000001010000011110011100110110;
   assign mem[11637] = 32'b11111011000010011101011101000000;
   assign mem[11638] = 32'b00000010000101010111100111011000;
   assign mem[11639] = 32'b11111111000111000001111110111100;
   assign mem[11640] = 32'b11111110001100101111011101111110;
   assign mem[11641] = 32'b00000100100001101011110101001000;
   assign mem[11642] = 32'b00001000010000100011100111010000;
   assign mem[11643] = 32'b11111011001011111101110011000000;
   assign mem[11644] = 32'b00001000000010100100110100000000;
   assign mem[11645] = 32'b11110111001101010000001100010000;
   assign mem[11646] = 32'b00000000000110000110101110111101;
   assign mem[11647] = 32'b00000100110011110000101100000000;
   assign mem[11648] = 32'b11110111100010110100010000000000;
   assign mem[11649] = 32'b11111001101100110000010110100000;
   assign mem[11650] = 32'b00000101101000100101000100110000;
   assign mem[11651] = 32'b11111010001011110110011001011000;
   assign mem[11652] = 32'b00000110011111010110111000101000;
   assign mem[11653] = 32'b00000110111001100010011100001000;
   assign mem[11654] = 32'b11110011111110100111110100100000;
   assign mem[11655] = 32'b00000011000000001110100010100000;
   assign mem[11656] = 32'b00000100010101101110000000011000;
   assign mem[11657] = 32'b00000000100001000000101000010110;
   assign mem[11658] = 32'b00000000001110110111111111011000;
   assign mem[11659] = 32'b11100100100000110111011111100000;
   assign mem[11660] = 32'b11110011011110000101101001110000;
   assign mem[11661] = 32'b00000100010001110001110101111000;
   assign mem[11662] = 32'b00000011101011101111110110110100;
   assign mem[11663] = 32'b00000010000100011111010001101000;
   assign mem[11664] = 32'b00000001010011000001101111000000;
   assign mem[11665] = 32'b11111011100010001011111100010000;
   assign mem[11666] = 32'b00000100010010001100001101000000;
   assign mem[11667] = 32'b11111110000010011101000001000000;
   assign mem[11668] = 32'b00000110101100111110001010101000;
   assign mem[11669] = 32'b11110111110110010110100111000000;
   assign mem[11670] = 32'b00000001000000010000010111010100;
   assign mem[11671] = 32'b11110100010101001100000000110000;
   assign mem[11672] = 32'b00000010001001001110010101101100;
   assign mem[11673] = 32'b00000010111000110000100110111100;
   assign mem[11674] = 32'b11111010100001101101100111100000;
   assign mem[11675] = 32'b00000100000010111001101111001000;
   assign mem[11676] = 32'b11111111111000101100101110010101;
   assign mem[11677] = 32'b00000000101100111101100010100000;
   assign mem[11678] = 32'b00000000000010000101100101011010;
   assign mem[11679] = 32'b11111011000001000100010000011000;
   assign mem[11680] = 32'b00000010101010111110001111010100;
   assign mem[11681] = 32'b00000011101011111000110111000100;
   assign mem[11682] = 32'b11111001010010100111100111010000;
   assign mem[11683] = 32'b11111100001011011111010011111000;
   assign mem[11684] = 32'b00000100110011101011011100110000;
   assign mem[11685] = 32'b11110110011111101101010101110000;
   assign mem[11686] = 32'b00001001111111110011000010110000;
   assign mem[11687] = 32'b11111111110011111111100100101111;
   assign mem[11688] = 32'b11111101010011000010110001110000;
   assign mem[11689] = 32'b00000011001001100100001101110000;
   assign mem[11690] = 32'b11110101100101001000011010010000;
   assign mem[11691] = 32'b11111000101101110010010011100000;
   assign mem[11692] = 32'b11110110001110000010111011000000;
   assign mem[11693] = 32'b00000010000101010011011011001000;
   assign mem[11694] = 32'b00001000101111111000110011100000;
   assign mem[11695] = 32'b11111100001010101101101110010000;
   assign mem[11696] = 32'b00000001101001011101110001110110;
   assign mem[11697] = 32'b00000101111101000001110010110000;
   assign mem[11698] = 32'b11111001010000101110011001111000;
   assign mem[11699] = 32'b00000111110110000100100000000000;
   assign mem[11700] = 32'b11110110011010101100001101110000;
   assign mem[11701] = 32'b11111111011010010001100011010100;
   assign mem[11702] = 32'b11111101010011010100011000001000;
   assign mem[11703] = 32'b00001000110000001010010100000000;
   assign mem[11704] = 32'b11111100011011010100101110010000;
   assign mem[11705] = 32'b00000001110011011001010011000100;
   assign mem[11706] = 32'b00000001101001001010110010111100;
   assign mem[11707] = 32'b11111010110111100000111110001000;
   assign mem[11708] = 32'b00001011001010111100101000100000;
   assign mem[11709] = 32'b11110010001110010110011001100000;
   assign mem[11710] = 32'b11111011010001010010101000101000;
   assign mem[11711] = 32'b11110111110111100111000000100000;
   assign mem[11712] = 32'b00000010101101110000100010010000;
   assign mem[11713] = 32'b00000100001000101010001010100000;
   assign mem[11714] = 32'b11111110111010000100101001100000;
   assign mem[11715] = 32'b11111111110000010000001110101000;
   assign mem[11716] = 32'b00000001010011011101111010000100;
   assign mem[11717] = 32'b11111000101101010111010100011000;
   assign mem[11718] = 32'b00000011001111000111100100001100;
   assign mem[11719] = 32'b11111101111101000101011111011000;
   assign mem[11720] = 32'b00000010100011100100011000110000;
   assign mem[11721] = 32'b11111110000110010000010100001010;
   assign mem[11722] = 32'b00000000110100110000010001011010;
   assign mem[11723] = 32'b11111101101010111110101111000100;
   assign mem[11724] = 32'b00000010101110011010001101100100;
   assign mem[11725] = 32'b11111011000011011100001001000000;
   assign mem[11726] = 32'b11111100001100101110100110111100;
   assign mem[11727] = 32'b00000011010001000100101000100000;
   assign mem[11728] = 32'b11110111100010101000010110110000;
   assign mem[11729] = 32'b00000001111110011111101110011010;
   assign mem[11730] = 32'b00000011001000000010100110011000;
   assign mem[11731] = 32'b00000011000000001100011010011100;
   assign mem[11732] = 32'b00000001110101101000011111000000;
   assign mem[11733] = 32'b11111111100100101100000010101010;
   assign mem[11734] = 32'b00000010100010001111111011100000;
   assign mem[11735] = 32'b00000010111010000000100000101000;
   assign mem[11736] = 32'b00000001100010010011001000011110;
   assign mem[11737] = 32'b11111101010001111001001000101100;
   assign mem[11738] = 32'b00000000111110010100101001001000;
   assign mem[11739] = 32'b11111101111111010001100111100000;
   assign mem[11740] = 32'b00000110001100000000100101011000;
   assign mem[11741] = 32'b11101111100101010011100010000000;
   assign mem[11742] = 32'b00000101010010000100101000100000;
   assign mem[11743] = 32'b00000100100011111100101000111000;
   assign mem[11744] = 32'b00000001101010100000111011110000;
   assign mem[11745] = 32'b11111110101000000101001100000000;
   assign mem[11746] = 32'b00000011110011111100100111111000;
   assign mem[11747] = 32'b11111111001111111000011010001100;
   assign mem[11748] = 32'b00000000110101000000111001100010;
   assign mem[11749] = 32'b00000010010101101000100010100100;
   assign mem[11750] = 32'b11111010110000101001011011000000;
   assign mem[11751] = 32'b00001000110111010001000100100000;
   assign mem[11752] = 32'b00000000011101111010010110000101;
   assign mem[11753] = 32'b00000001001100001011111000110010;
   assign mem[11754] = 32'b11111101100100010001011010110100;
   assign mem[11755] = 32'b00000000111100001001110011111010;
   assign mem[11756] = 32'b11111111010000010111101101100111;
   assign mem[11757] = 32'b11111001001001001101010000101000;
   assign mem[11758] = 32'b11111111110101100000101000000001;
   assign mem[11759] = 32'b00000000110100101001001100111010;
   assign mem[11760] = 32'b00000000110100111000110111000000;
   assign mem[11761] = 32'b00000011001010011001101101101100;
   assign mem[11762] = 32'b11111000000000001011101000001000;
   assign mem[11763] = 32'b00000010000001011110111011011000;
   assign mem[11764] = 32'b11111111010011001100000001101000;
   assign mem[11765] = 32'b00000010000011111000001101000100;
   assign mem[11766] = 32'b00000001000101011101010111001100;
   assign mem[11767] = 32'b11111110100110101001011011010110;
   assign mem[11768] = 32'b00000001101111000011011111010010;
   assign mem[11769] = 32'b00000000110110001000100110100111;
   assign mem[11770] = 32'b11111011010111101110101011010000;
   assign mem[11771] = 32'b00000010011011011110010000100000;
   assign mem[11772] = 32'b00000000110000111010011101001100;
   assign mem[11773] = 32'b00000000011000110100100000100100;
   assign mem[11774] = 32'b00000001010100101101001010111110;
   assign mem[11775] = 32'b00000010000010101111011101000100;
   assign mem[11776] = 32'b11111101001100111101001100010000;
   assign mem[11777] = 32'b00000001010000110001010011100110;
   assign mem[11778] = 32'b00000001111010100000110100101110;
   assign mem[11779] = 32'b00000010101100101111011101101100;
   assign mem[11780] = 32'b11111101100111000101011011001100;
   assign mem[11781] = 32'b00000001100110010101010000111110;
   assign mem[11782] = 32'b11111100111110010001111110000100;
   assign mem[11783] = 32'b11111101110010110001001111001100;
   assign mem[11784] = 32'b11111110000100000010111011010110;
   assign mem[11785] = 32'b11111010000111010010101011010000;
   assign mem[11786] = 32'b11111111001110010111101100101011;
   assign mem[11787] = 32'b11111110100001010010001101001000;
   assign mem[11788] = 32'b00000010100000111001011000111000;
   assign mem[11789] = 32'b11111111001000110111111011011010;
   assign mem[11790] = 32'b00000101010110111010100101000000;
   assign mem[11791] = 32'b00010010011011110110010100100000;
   assign mem[11792] = 32'b00001110000001111011010011110000;
   assign mem[11793] = 32'b11110011111001001101001100110000;
   assign mem[11794] = 32'b11110111001000011001010001000000;
   assign mem[11795] = 32'b00000010101010011110001001000100;
   assign mem[11796] = 32'b11110001110111010011000001110000;
   assign mem[11797] = 32'b00001001101110010001111010010000;
   assign mem[11798] = 32'b11101110100001010011010101100000;
   assign mem[11799] = 32'b00000010000110010010100010011000;
   assign mem[11800] = 32'b11111011100001001001100101001000;
   assign mem[11801] = 32'b11111101011111110010000100100000;
   assign mem[11802] = 32'b00000001000001110001111100101100;
   assign mem[11803] = 32'b11111111111100100001111110111101;
   assign mem[11804] = 32'b00000101001111000111110110100000;
   assign mem[11805] = 32'b11111011111111111100101011001000;
   assign mem[11806] = 32'b00000101111111101111101101010000;
   assign mem[11807] = 32'b00000001101110010000101111110000;
   assign mem[11808] = 32'b00000000011011111010100010010000;
   assign mem[11809] = 32'b11110100010100011110100100010000;
   assign mem[11810] = 32'b00001001010110111110100110010000;
   assign mem[11811] = 32'b11110011100110000010011111000000;
   assign mem[11812] = 32'b00000110110001000110011101010000;
   assign mem[11813] = 32'b11111011100011111011110001001000;
   assign mem[11814] = 32'b11110111110010001100110110000000;
   assign mem[11815] = 32'b00000001001010110110010110100100;
   assign mem[11816] = 32'b00000100000110110101011100111000;
   assign mem[11817] = 32'b11110011111101110001100000110000;
   assign mem[11818] = 32'b11101111001101010111100000000000;
   assign mem[11819] = 32'b11111101111010101011101100100000;
   assign mem[11820] = 32'b00000010011000010101101011001100;
   assign mem[11821] = 32'b00000001101110001001111010011100;
   assign mem[11822] = 32'b11111110010100001101010111010000;
   assign mem[11823] = 32'b00000000000110010111010001110011;
   assign mem[11824] = 32'b00000001000000111010100100010010;
   assign mem[11825] = 32'b00000000110100100001011100010011;
   assign mem[11826] = 32'b11111011110010010111001000110000;
   assign mem[11827] = 32'b00000010010101101010010010010000;
   assign mem[11828] = 32'b11111100001011100010011111000000;
   assign mem[11829] = 32'b00000010110001011000100100101100;
   assign mem[11830] = 32'b00000011100000100101001100001100;
   assign mem[11831] = 32'b11111011110001000010111100010000;
   assign mem[11832] = 32'b11111110000110110010110010010000;
   assign mem[11833] = 32'b11111100101011111000011111111100;
   assign mem[11834] = 32'b00000100001111000010101000111000;
   assign mem[11835] = 32'b11111110000001000110110110011110;
   assign mem[11836] = 32'b00000011011100001010011010011100;
   assign mem[11837] = 32'b00000110011001100000011000100000;
   assign mem[11838] = 32'b11111111101111110101101001000001;
   assign mem[11839] = 32'b11110111111101100100010111010000;
   assign mem[11840] = 32'b11111100100000001100011110111000;
   assign mem[11841] = 32'b11111010011101001100001011000000;
   assign mem[11842] = 32'b00000100110011111010010001000000;
   assign mem[11843] = 32'b00000110111000010001011001101000;
   assign mem[11844] = 32'b11111110011110101110010101100010;
   assign mem[11845] = 32'b11111101101111111001000001110000;
   assign mem[11846] = 32'b00000100010101010101000010100000;
   assign mem[11847] = 32'b11111111110011010110001101110110;
   assign mem[11848] = 32'b11111101011010101101010100011000;
   assign mem[11849] = 32'b11111011100011110111110110010000;
   assign mem[11850] = 32'b00001000111001000101101110100000;
   assign mem[11851] = 32'b00000000100010011100010011110111;
   assign mem[11852] = 32'b00001000110011110101100110100000;
   assign mem[11853] = 32'b11110111011101011010100100010000;
   assign mem[11854] = 32'b00000000001100101110111100000100;
   assign mem[11855] = 32'b00000011010011111101100101110000;
   assign mem[11856] = 32'b00000100011111001001011000100000;
   assign mem[11857] = 32'b00000001011110100010000001100000;
   assign mem[11858] = 32'b11111010110100111110001110100000;
   assign mem[11859] = 32'b11111100011011101111001111001100;
   assign mem[11860] = 32'b11111010110010111111111100101000;
   assign mem[11861] = 32'b11111111000011011111010011100101;
   assign mem[11862] = 32'b00000000000111011010110010011101;
   assign mem[11863] = 32'b00000000000100111110011100010000;
   assign mem[11864] = 32'b00000101001011010100000001111000;
   assign mem[11865] = 32'b11111010000010110011010000111000;
   assign mem[11866] = 32'b00000000111100011101011001110110;
   assign mem[11867] = 32'b00000110010000110111001101111000;
   assign mem[11868] = 32'b00000001011011101100001000000010;
   assign mem[11869] = 32'b11111010111011100100011001110000;
   assign mem[11870] = 32'b00000001000011100101001011100110;
   assign mem[11871] = 32'b00000011100000111010101111110100;
   assign mem[11872] = 32'b00000000011000110101110000011101;
   assign mem[11873] = 32'b11111110010011100000110100100010;
   assign mem[11874] = 32'b11111100100100110111100110001100;
   assign mem[11875] = 32'b00000001110110000110101011111000;
   assign mem[11876] = 32'b11111101110111101100101110011000;
   assign mem[11877] = 32'b00000011001100000011001010101100;
   assign mem[11878] = 32'b11110101110110011101111001110000;
   assign mem[11879] = 32'b00000011101100101011111110110100;
   assign mem[11880] = 32'b00000000001101110100000001011011;
   assign mem[11881] = 32'b11110111010000111111011000010000;
   assign mem[11882] = 32'b00000001110110101110001000010010;
   assign mem[11883] = 32'b00001000111011000000100101010000;
   assign mem[11884] = 32'b11110010011010000011010001000000;
   assign mem[11885] = 32'b00000110000010111101101010001000;
   assign mem[11886] = 32'b00000001011001001100110110000010;
   assign mem[11887] = 32'b11111011110101100000110001111000;
   assign mem[11888] = 32'b00001001111111011000111100110000;
   assign mem[11889] = 32'b11100001000110101001110110100000;
   assign mem[11890] = 32'b11111100010110111010110101001100;
   assign mem[11891] = 32'b11111011000011101111101100110000;
   assign mem[11892] = 32'b00000010011001100111001111010100;
   assign mem[11893] = 32'b00000111110001100100111000000000;
   assign mem[11894] = 32'b11111010001011100111110110001000;
   assign mem[11895] = 32'b00000101010000111101001011100000;
   assign mem[11896] = 32'b00001001001000001110001110010000;
   assign mem[11897] = 32'b11111000010101101101010101100000;
   assign mem[11898] = 32'b00000101000111100001011000111000;
   assign mem[11899] = 32'b11101100011001111011111110000000;
   assign mem[11900] = 32'b11110111110111010010011101000000;
   assign mem[11901] = 32'b00000101000010110000010111110000;
   assign mem[11902] = 32'b11111101001000100111110110010000;
   assign mem[11903] = 32'b11111001110111110001101110101000;
   assign mem[11904] = 32'b00001010011000111101011001010000;
   assign mem[11905] = 32'b11111101110010111011011001000100;
   assign mem[11906] = 32'b00000110110110101100011111011000;
   assign mem[11907] = 32'b00000101000001100111010110101000;
   assign mem[11908] = 32'b11111100010010000110010001110100;
   assign mem[11909] = 32'b00000010101000010111010011111100;
   assign mem[11910] = 32'b11111011010011000010011101010000;
   assign mem[11911] = 32'b11110101110100010100000111010000;
   assign mem[11912] = 32'b00000011000111111010111000010100;
   assign mem[11913] = 32'b00000000000000011110011110010000;
   assign mem[11914] = 32'b11110011100000111110101001000000;
   assign mem[11915] = 32'b11111110111100001000011100010000;
   assign mem[11916] = 32'b11111000101011010111101110001000;
   assign mem[11917] = 32'b00000110101100101011100011101000;
   assign mem[11918] = 32'b00000011110110001010110000101000;
   assign mem[11919] = 32'b00000100100011111111001110011000;
   assign mem[11920] = 32'b11111000111010100110000010010000;
   assign mem[11921] = 32'b11111100010011111010110011101000;
   assign mem[11922] = 32'b00000000100010110000000110110100;
   assign mem[11923] = 32'b11111101110110000011010111010000;
   assign mem[11924] = 32'b00000100010011100110101010010000;
   assign mem[11925] = 32'b00000100011110001111101110110000;
   assign mem[11926] = 32'b00000010100110100110000010010000;
   assign mem[11927] = 32'b11111101110000011101000110010000;
   assign mem[11928] = 32'b00000010101100011100011111110100;
   assign mem[11929] = 32'b00000011110110000010111001100000;
   assign mem[11930] = 32'b00000001110100111100100111101100;
   assign mem[11931] = 32'b00001001011100101110000111010000;
   assign mem[11932] = 32'b11111110000000110110001101111100;
   assign mem[11933] = 32'b11111000101110111110011010111000;
   assign mem[11934] = 32'b00000111010001110110111100010000;
   assign mem[11935] = 32'b11110100101101100011110101010000;
   assign mem[11936] = 32'b11111111001010101101100100001010;
   assign mem[11937] = 32'b00000011011100001101110111000100;
   assign mem[11938] = 32'b11111111010000010100010010100001;
   assign mem[11939] = 32'b00001000110101100101110001010000;
   assign mem[11940] = 32'b11111111101110011011010000000001;
   assign mem[11941] = 32'b00001011101010101110101101110000;
   assign mem[11942] = 32'b11111111001110000010110111111001;
   assign mem[11943] = 32'b00000010111110101011100010110000;
   assign mem[11944] = 32'b11111001001000101011001011010000;
   assign mem[11945] = 32'b00000010011010001110110101010000;
   assign mem[11946] = 32'b00000000000000100001010011011100;
   assign mem[11947] = 32'b11111001100110111110110011001000;
   assign mem[11948] = 32'b00000001100000001100101101100110;
   assign mem[11949] = 32'b11110110100100111011110111100000;
   assign mem[11950] = 32'b11111001000000110011010110101000;
   assign mem[11951] = 32'b11111111101111010011100000110111;
   assign mem[11952] = 32'b11111100101001000100011101101100;
   assign mem[11953] = 32'b00000100000100100010101110110000;
   assign mem[11954] = 32'b11111001111000110011011110111000;
   assign mem[11955] = 32'b00000011110010100111000001001100;
   assign mem[11956] = 32'b00000011111100001111111110010000;
   assign mem[11957] = 32'b11111011000110001110111100110000;
   assign mem[11958] = 32'b00000010101111110100110101000000;
   assign mem[11959] = 32'b00000000011110010011111101110111;
   assign mem[11960] = 32'b11111011100001010011010010010000;
   assign mem[11961] = 32'b00001010100001100010110100100000;
   assign mem[11962] = 32'b11111100010100001110010010001100;
   assign mem[11963] = 32'b11111101100110010111000011110100;
   assign mem[11964] = 32'b00000111100010111111111101101000;
   assign mem[11965] = 32'b11111110111001011110011101011110;
   assign mem[11966] = 32'b00000110110001000010010100011000;
   assign mem[11967] = 32'b00000110000110001101101100011000;
   assign mem[11968] = 32'b11111010011000110000000000011000;
   assign mem[11969] = 32'b11111000001111110111001101010000;
   assign mem[11970] = 32'b11110001110100010100110011100000;
   assign mem[11971] = 32'b11110111100001010100011100110000;
   assign mem[11972] = 32'b00001001011110000111000000000000;
   assign mem[11973] = 32'b00000101010011010001110001101000;
   assign mem[11974] = 32'b00000100100011101101101011001000;
   assign mem[11975] = 32'b00001000010010011010001101000000;
   assign mem[11976] = 32'b00000101010101000010001111110000;
   assign mem[11977] = 32'b11110010101010010111011100110000;
   assign mem[11978] = 32'b00000001010100011111100011011000;
   assign mem[11979] = 32'b11111000100101001001100110110000;
   assign mem[11980] = 32'b00000000101100111011001111111001;
   assign mem[11981] = 32'b11110101101100111011000111000000;
   assign mem[11982] = 32'b00000000001001111111001111110111;
   assign mem[11983] = 32'b11111101100111100010001000100100;
   assign mem[11984] = 32'b00000001010100101111101011101000;
   assign mem[11985] = 32'b11111111000111000111101000010111;
   assign mem[11986] = 32'b11111100011001010110110111110100;
   assign mem[11987] = 32'b00000010010111011110101000010000;
   assign mem[11988] = 32'b11111100000101111011000100000100;
   assign mem[11989] = 32'b00000101101100010101101110001000;
   assign mem[11990] = 32'b11111110011000110110111001101110;
   assign mem[11991] = 32'b11111111111101001101110101011010;
   assign mem[11992] = 32'b11111100101100100000100101010100;
   assign mem[11993] = 32'b11111011101011101011111111100000;
   assign mem[11994] = 32'b00000010010101011110110010111000;
   assign mem[11995] = 32'b11111101100110110000100101010100;
   assign mem[11996] = 32'b11111011101100100100111100100000;
   assign mem[11997] = 32'b00000010100110101000101010111000;
   assign mem[11998] = 32'b00000000101010100010110111100011;
   assign mem[11999] = 32'b11111101001000100010010000100000;
   assign mem[12000] = 32'b11111011001010100101010100010000;
   assign mem[12001] = 32'b00000010110101011010111111001000;
   assign mem[12002] = 32'b00000000001010111111010110100011;
   assign mem[12003] = 32'b11111100110001101101110010000000;
   assign mem[12004] = 32'b00000100111010001000001111110000;
   assign mem[12005] = 32'b11111010101110101010000011011000;
   assign mem[12006] = 32'b11111111100010010010100000110001;
   assign mem[12007] = 32'b00000011010010000000010110011100;
   assign mem[12008] = 32'b11111101000010100011011011001100;
   assign mem[12009] = 32'b11111111000000111111000101001001;
   assign mem[12010] = 32'b00000001110001010000011011011010;
   assign mem[12011] = 32'b11110111111001111101011001010000;
   assign mem[12012] = 32'b00001000010100010001111001110000;
   assign mem[12013] = 32'b11111111100110110101110100011010;
   assign mem[12014] = 32'b00000011001000100011110111110000;
   assign mem[12015] = 32'b11111100010001001011010100010000;
   assign mem[12016] = 32'b11111100011110101111011010100100;
   assign mem[12017] = 32'b00001001111000011110010010010000;
   assign mem[12018] = 32'b11110111010110111011010010100000;
   assign mem[12019] = 32'b00000001111101000100101101000000;
   assign mem[12020] = 32'b11111111110110100011101001100000;
   assign mem[12021] = 32'b11110011100101110000111101010000;
   assign mem[12022] = 32'b00000001111100011010010011010000;
   assign mem[12023] = 32'b00000011001011010011101100001100;
   assign mem[12024] = 32'b11111010111010010110010010011000;
   assign mem[12025] = 32'b00000010001010000010101100111100;
   assign mem[12026] = 32'b00000010001110100001111110001000;
   assign mem[12027] = 32'b11110111011101110101111011110000;
   assign mem[12028] = 32'b00000011001000110100101110001000;
   assign mem[12029] = 32'b11111111101111101110010110110111;
   assign mem[12030] = 32'b00000110011011011100010111010000;
   assign mem[12031] = 32'b00000100101101010000001100110000;
   assign mem[12032] = 32'b11110001101010010110011011000000;
   assign mem[12033] = 32'b11111011111101110100110011001000;
   assign mem[12034] = 32'b00000001101000100000010010111110;
   assign mem[12035] = 32'b00000011011001110001110101111000;
   assign mem[12036] = 32'b11111111111110011100111001111110;
   assign mem[12037] = 32'b00001010110000111001011000100000;
   assign mem[12038] = 32'b11110100101110000101101101110000;
   assign mem[12039] = 32'b00000010011100110001000011111100;
   assign mem[12040] = 32'b00000011101000000000011100101000;
   assign mem[12041] = 32'b11111010000100111111001100001000;
   assign mem[12042] = 32'b00000011110000010100001000001100;
   assign mem[12043] = 32'b11111111001011010101000100100110;
   assign mem[12044] = 32'b00000010111001000111001010101000;
   assign mem[12045] = 32'b11111101110000000011111011110000;
   assign mem[12046] = 32'b00000101110100010110011101101000;
   assign mem[12047] = 32'b11111110101000000101110011011100;
   assign mem[12048] = 32'b00000001010111001010011000000100;
   assign mem[12049] = 32'b11111001000110011010110010111000;
   assign mem[12050] = 32'b11111110111011010100110100010000;
   assign mem[12051] = 32'b11111011010100111011110111111000;
   assign mem[12052] = 32'b00000001110010101011110000010010;
   assign mem[12053] = 32'b00000101000011111100011011111000;
   assign mem[12054] = 32'b00000000110111100010001111000111;
   assign mem[12055] = 32'b00000010100000000111001010001000;
   assign mem[12056] = 32'b00000001011001101000111111111100;
   assign mem[12057] = 32'b00000011001101111101101111010000;
   assign mem[12058] = 32'b00000001100110101100110010111000;
   assign mem[12059] = 32'b11110011001100011100100111000000;
   assign mem[12060] = 32'b00000101010100000001101101010000;
   assign mem[12061] = 32'b11110110111011011000010101010000;
   assign mem[12062] = 32'b11111101100111101110110001110100;
   assign mem[12063] = 32'b00000001011110001100111111100010;
   assign mem[12064] = 32'b00000010001000100110101001000100;
   assign mem[12065] = 32'b11111111010101010001010101110011;
   assign mem[12066] = 32'b00000011000101100010000001000100;
   assign mem[12067] = 32'b00000100110001101101100111000000;
   assign mem[12068] = 32'b11111111011101011100001000101011;
   assign mem[12069] = 32'b00000010100000010101011011111100;
   assign mem[12070] = 32'b00000101111110110010110110110000;
   assign mem[12071] = 32'b00000100101010111010111101000000;
   assign mem[12072] = 32'b00000010011000111001010110101000;
   assign mem[12073] = 32'b11111110001011100110100101000100;
   assign mem[12074] = 32'b11111011001000100001111010111000;
   assign mem[12075] = 32'b00000000001001010000100100000011;
   assign mem[12076] = 32'b11111110000111101011010010101100;
   assign mem[12077] = 32'b00000001111001100010001110110110;
   assign mem[12078] = 32'b11111011100001001100000010010000;
   assign mem[12079] = 32'b00000000000110000110101100000010;
   assign mem[12080] = 32'b00000001010000001110110111101110;
   assign mem[12081] = 32'b11111111000001100111111100011111;
   assign mem[12082] = 32'b11111011101001111001100111101000;
   assign mem[12083] = 32'b00000100011111001011010111000000;
   assign mem[12084] = 32'b11111011110010010010001100110000;
   assign mem[12085] = 32'b00000001000011010010110011010100;
   assign mem[12086] = 32'b00001001110100001111101111010000;
   assign mem[12087] = 32'b11111100100000001000110100101100;
   assign mem[12088] = 32'b11111101111111111010010010110000;
   assign mem[12089] = 32'b00000101100011111100100001010000;
   assign mem[12090] = 32'b11111000011000011000100101011000;
   assign mem[12091] = 32'b00000011111111100111010111100000;
   assign mem[12092] = 32'b11111101001101001011110111011100;
   assign mem[12093] = 32'b00000110011100011101011100101000;
   assign mem[12094] = 32'b11111110100010000010100110000110;
   assign mem[12095] = 32'b00000110000011101101100100100000;
   assign mem[12096] = 32'b11111111111101110011000001100100;
   assign mem[12097] = 32'b11111100101001110100100011100000;
   assign mem[12098] = 32'b00000011010110110110100000111100;
   assign mem[12099] = 32'b11111101010011001011101101000000;
   assign mem[12100] = 32'b00001001100000010100000010100000;
   assign mem[12101] = 32'b00000001000000111101110011000100;
   assign mem[12102] = 32'b11111111000000111101100011100001;
   assign mem[12103] = 32'b11111010110100100000111101101000;
   assign mem[12104] = 32'b11101101100000001001110010100000;
   assign mem[12105] = 32'b00000100111000011110100111001000;
   assign mem[12106] = 32'b00000011011100011011110000101000;
   assign mem[12107] = 32'b11111110110010101011011011000000;
   assign mem[12108] = 32'b11111000101100001000001011001000;
   assign mem[12109] = 32'b11110100111100101101010001100000;
   assign mem[12110] = 32'b11111111011001001111010000000010;
   assign mem[12111] = 32'b11111111111101000000010111110010;
   assign mem[12112] = 32'b00000001111010011010110011010000;
   assign mem[12113] = 32'b00000000000101110110100001101100;
   assign mem[12114] = 32'b11111100000000111010101011010000;
   assign mem[12115] = 32'b00000011100000100010101011110100;
   assign mem[12116] = 32'b00000011000010010010100000100000;
   assign mem[12117] = 32'b11111010001111100000100110101000;
   assign mem[12118] = 32'b00000001110000111000101000110100;
   assign mem[12119] = 32'b11111000111011000110101001110000;
   assign mem[12120] = 32'b00000001000010111100111001011100;
   assign mem[12121] = 32'b11110100000110001111000110100000;
   assign mem[12122] = 32'b00001010111001010100100011010000;
   assign mem[12123] = 32'b00000010011010010010111100011000;
   assign mem[12124] = 32'b11110101110110110110111110000000;
   assign mem[12125] = 32'b11111111000010110110111100101011;
   assign mem[12126] = 32'b11111100101100110011011000010000;
   assign mem[12127] = 32'b00001001001000110010001110110000;
   assign mem[12128] = 32'b00000010000010100110010100001000;
   assign mem[12129] = 32'b00000011011111011001110111100000;
   assign mem[12130] = 32'b00000100010110110100100001001000;
   assign mem[12131] = 32'b11111000010001111111011111010000;
   assign mem[12132] = 32'b00000011100111100110101001011000;
   assign mem[12133] = 32'b11111010010011111010011000110000;
   assign mem[12134] = 32'b11111100100101001010000000101000;
   assign mem[12135] = 32'b11111111100001011001100111010100;
   assign mem[12136] = 32'b00000000101100110001110001100011;
   assign mem[12137] = 32'b00000111011110010110011101111000;
   assign mem[12138] = 32'b11111000101011011110001101011000;
   assign mem[12139] = 32'b11111101000111111100110001000000;
   assign mem[12140] = 32'b00000010110110111001101011010000;
   assign mem[12141] = 32'b00001000111110111001011001000000;
   assign mem[12142] = 32'b00000001100111010010001011101000;
   assign mem[12143] = 32'b11110100011110111110111001000000;
   assign mem[12144] = 32'b11111110101110100110001110101110;
   assign mem[12145] = 32'b11111010000001010100001001000000;
   assign mem[12146] = 32'b11110111100011101000110011000000;
   assign mem[12147] = 32'b00001010011101001011011101100000;
   assign mem[12148] = 32'b11110001111010100000111000110000;
   assign mem[12149] = 32'b00000001011000000101001101110010;
   assign mem[12150] = 32'b00000010010001101111011011001100;
   assign mem[12151] = 32'b00000010000001101010110110101000;
   assign mem[12152] = 32'b00000010001011010111111100111000;
   assign mem[12153] = 32'b00000001011001011001100111111100;
   assign mem[12154] = 32'b11111101110110110001001100110100;
   assign mem[12155] = 32'b11111100101010011110001100010000;
   assign mem[12156] = 32'b11111101111101010101000111011100;
   assign mem[12157] = 32'b00000011001011011010110100010000;
   assign mem[12158] = 32'b11111001000110110100110010100000;
   assign mem[12159] = 32'b11111111100000100011101111001001;
   assign mem[12160] = 32'b00000001111111101011110110011000;
   assign mem[12161] = 32'b00000010010100011100011101101100;
   assign mem[12162] = 32'b00000101010110110011111001100000;
   assign mem[12163] = 32'b11111101001011110111100000011100;
   assign mem[12164] = 32'b11110100000001100110010010010000;
   assign mem[12165] = 32'b11110110101000010101111000100000;
   assign mem[12166] = 32'b00000001100011101110000010110010;
   assign mem[12167] = 32'b00000101000000001100011001010000;
   assign mem[12168] = 32'b11111100000110110001000111100000;
   assign mem[12169] = 32'b11111101101000000101011101111100;
   assign mem[12170] = 32'b11111001111000100100000000011000;
   assign mem[12171] = 32'b11111101011000011010011010010000;
   assign mem[12172] = 32'b11111100110011000010011100000000;
   assign mem[12173] = 32'b00000100000111111010110010000000;
   assign mem[12174] = 32'b11110111111011101010000000010000;
   assign mem[12175] = 32'b00000010110011011000001100110100;
   assign mem[12176] = 32'b00001000111110100011100101000000;
   assign mem[12177] = 32'b11111001001100001101010111000000;
   assign mem[12178] = 32'b00000100000000001101000011000000;
   assign mem[12179] = 32'b11111011001101101101111001001000;
   assign mem[12180] = 32'b11111011000010110101100110111000;
   assign mem[12181] = 32'b11111011100001110000000111001000;
   assign mem[12182] = 32'b00000011110000100110111111100100;
   assign mem[12183] = 32'b00000000111000111001011111001000;
   assign mem[12184] = 32'b11111101010111111000101000100000;
   assign mem[12185] = 32'b00000100001111111100010111010000;
   assign mem[12186] = 32'b00000010101011100010010010001100;
   assign mem[12187] = 32'b11111000110010001000011100101000;
   assign mem[12188] = 32'b00000101001000000001101100110000;
   assign mem[12189] = 32'b00000000000110111011000101001101;
   assign mem[12190] = 32'b00000000111000100110100001010011;
   assign mem[12191] = 32'b11111010101000011100010001001000;
   assign mem[12192] = 32'b00001101010010101010000101000000;
   assign mem[12193] = 32'b11110110001111001111010000000000;
   assign mem[12194] = 32'b00000100101110001110010010110000;
   assign mem[12195] = 32'b11111010100000011011010011000000;
   assign mem[12196] = 32'b11111011101001011110011001000000;
   assign mem[12197] = 32'b00000110110001010011101101000000;
   assign mem[12198] = 32'b11111110111110111100001111110100;
   assign mem[12199] = 32'b11101100111011000000101110000000;
   assign mem[12200] = 32'b00001011110101011101001010010000;
   assign mem[12201] = 32'b00000000001001110111111001011111;
   assign mem[12202] = 32'b00001010111111000110101011100000;
   assign mem[12203] = 32'b11101011000000100000011000000000;
   assign mem[12204] = 32'b00000100000010111100011100000000;
   assign mem[12205] = 32'b11110111110000100110101100100000;
   assign mem[12206] = 32'b11111011000000011100110011100000;
   assign mem[12207] = 32'b11111111110101001011111110101000;
   assign mem[12208] = 32'b00000010110001000011110101100000;
   assign mem[12209] = 32'b11111010110011110001100110101000;
   assign mem[12210] = 32'b00000011001010011011001011110000;
   assign mem[12211] = 32'b11111010100101101101001011001000;
   assign mem[12212] = 32'b00000010111011001010011000110100;
   assign mem[12213] = 32'b00000000001001001101001100100011;
   assign mem[12214] = 32'b00000001011011101000011001010000;
   assign mem[12215] = 32'b11111101000000100011010001010000;
   assign mem[12216] = 32'b00000000001101011011101011111100;
   assign mem[12217] = 32'b00000101110000100100010011111000;
   assign mem[12218] = 32'b11110010000010101101100100010000;
   assign mem[12219] = 32'b11111110111111000110000011001100;
   assign mem[12220] = 32'b00000100000000000110000001110000;
   assign mem[12221] = 32'b11111101100000000000011101100000;
   assign mem[12222] = 32'b11111111010101001110010000110001;
   assign mem[12223] = 32'b00000010000001111011110010000000;
   assign mem[12224] = 32'b00000001000001110110000010010100;
   assign mem[12225] = 32'b11111101000111100001101000111100;
   assign mem[12226] = 32'b11111111110011100010000001101110;
   assign mem[12227] = 32'b00000001110011001100011101001010;
   assign mem[12228] = 32'b00000001110001100100110011110110;
   assign mem[12229] = 32'b00000001111011011100010011110110;
   assign mem[12230] = 32'b00000101110001111110010111001000;
   assign mem[12231] = 32'b11111110110100010100110101011000;
   assign mem[12232] = 32'b00000001110000000110001010000000;
   assign mem[12233] = 32'b11111010100101111110111010111000;
   assign mem[12234] = 32'b11111010000011101111000010110000;
   assign mem[12235] = 32'b11110101100011011011000010000000;
   assign mem[12236] = 32'b00000101101110110001000101110000;
   assign mem[12237] = 32'b00000010000101110010111001110000;
   assign mem[12238] = 32'b00000000001111110010000001101001;
   assign mem[12239] = 32'b11111110110000111010111101110000;
   assign mem[12240] = 32'b11110111100111001100100100100000;
   assign mem[12241] = 32'b00000101001011111010110010000000;
   assign mem[12242] = 32'b00000100010100011111000101001000;
   assign mem[12243] = 32'b11110111111111101101001100110000;
   assign mem[12244] = 32'b11111111101110000011000100010101;
   assign mem[12245] = 32'b00000110000000101011010001011000;
   assign mem[12246] = 32'b11111111101000101101111100110110;
   assign mem[12247] = 32'b00000110000010110100001011101000;
   assign mem[12248] = 32'b00000000010001001111001001011110;
   assign mem[12249] = 32'b11110010101111001000010010000000;
   assign mem[12250] = 32'b00000010111100001101011001010000;
   assign mem[12251] = 32'b11111101111110110110110111100000;
   assign mem[12252] = 32'b11110001010010010110111000000000;
   assign mem[12253] = 32'b00000000111001100111001010010001;
   assign mem[12254] = 32'b00000000010001110010111001101101;
   assign mem[12255] = 32'b11110110111010110100001000100000;
   assign mem[12256] = 32'b00001011010010000001101100010000;
   assign mem[12257] = 32'b00000011000101001001011111001000;
   assign mem[12258] = 32'b11111000000000001011001001101000;
   assign mem[12259] = 32'b00000110110000110111000110010000;
   assign mem[12260] = 32'b00000001010110111000000101011110;
   assign mem[12261] = 32'b00000001111011110000011101110000;
   assign mem[12262] = 32'b00000110001101101111100101011000;
   assign mem[12263] = 32'b11110001011111011110011000100000;
   assign mem[12264] = 32'b00001001001101001010010111110000;
   assign mem[12265] = 32'b11110111100100100010100100010000;
   assign mem[12266] = 32'b11110011101011010010001011110000;
   assign mem[12267] = 32'b00000101001000110100111101000000;
   assign mem[12268] = 32'b11110100010111001001010011110000;
   assign mem[12269] = 32'b11110101110011111110100101010000;
   assign mem[12270] = 32'b11111111010111111110001011111011;
   assign mem[12271] = 32'b11110100000001000101111101100000;
   assign mem[12272] = 32'b00000110011011000110110111001000;
   assign mem[12273] = 32'b00000000111000010110000100010010;
   assign mem[12274] = 32'b00000100100100010011001110011000;
   assign mem[12275] = 32'b11111101000111111101011000010000;
   assign mem[12276] = 32'b11111100011011001101111011111100;
   assign mem[12277] = 32'b11111000111110111010001110010000;
   assign mem[12278] = 32'b00000010010010111001110100000100;
   assign mem[12279] = 32'b11111011011010111111001000101000;
   assign mem[12280] = 32'b11101101111110000110100110100000;
   assign mem[12281] = 32'b00000110011111000100010000000000;
   assign mem[12282] = 32'b00001100111101000010110011000000;
   assign mem[12283] = 32'b11111000001001000100011000111000;
   assign mem[12284] = 32'b00001010100101000100110111100000;
   assign mem[12285] = 32'b11111011100011010110010101100000;
   assign mem[12286] = 32'b11111000011100111100101010010000;
   assign mem[12287] = 32'b00001010010100010010000010110000;
   assign mem[12288] = 32'b11110101000110010100111001100000;
   assign mem[12289] = 32'b00000000001001111011011100101011;
   assign mem[12290] = 32'b11100001100101011001110100100000;
   assign mem[12291] = 32'b00000011100100000101100010111000;
   assign mem[12292] = 32'b00000011010100011011010101101000;
   assign mem[12293] = 32'b11111110001101011000101100011100;
   assign mem[12294] = 32'b00000011110001000011011110000000;
   assign mem[12295] = 32'b11111101000000111011111000010100;
   assign mem[12296] = 32'b11111110110001011110110101111110;
   assign mem[12297] = 32'b00000110110100110010000000110000;
   assign mem[12298] = 32'b11111111000100101011000100111101;
   assign mem[12299] = 32'b11110111010111001010011010110000;
   assign mem[12300] = 32'b11110111101010101001101000110000;
   assign mem[12301] = 32'b00000000101101000111010111101110;
   assign mem[12302] = 32'b00000101011111110010000000110000;
   assign mem[12303] = 32'b00000010100101101111100001000000;
   assign mem[12304] = 32'b00000110011110010101110010100000;
   assign mem[12305] = 32'b11111101000101111011110101011100;
   assign mem[12306] = 32'b11111110000010011101000100111010;
   assign mem[12307] = 32'b00000100110110110110111100111000;
   assign mem[12308] = 32'b00000000111001010001010101000101;
   assign mem[12309] = 32'b00000001111111011010111000000000;
   assign mem[12310] = 32'b00000101001000010111010111000000;
   assign mem[12311] = 32'b11110111100011100001101001000000;
   assign mem[12312] = 32'b11110010110000001111101100000000;
   assign mem[12313] = 32'b11111100111100001001110010001100;
   assign mem[12314] = 32'b11111001100110011000110110110000;
   assign mem[12315] = 32'b11111100100010110001100010100100;
   assign mem[12316] = 32'b00000000111000001110100110010000;
   assign mem[12317] = 32'b00000110001001000110100101100000;
   assign mem[12318] = 32'b00000000001010000101100110100111;
   assign mem[12319] = 32'b11111001110110000000101010011000;
   assign mem[12320] = 32'b00000100001011110101000111100000;
   assign mem[12321] = 32'b11111011000010011111101001110000;
   assign mem[12322] = 32'b00000011101001110010010110011100;
   assign mem[12323] = 32'b11110111010100010110011000010000;
   assign mem[12324] = 32'b00000000111011001100011000111101;
   assign mem[12325] = 32'b11101111010011111100110010000000;
   assign mem[12326] = 32'b00001000001010100011001001100000;
   assign mem[12327] = 32'b00000101101000110100101111001000;
   assign mem[12328] = 32'b11111011100110011100001110000000;
   assign mem[12329] = 32'b11110100001010001111010101010000;
   assign mem[12330] = 32'b11111011111001000000111110101000;
   assign mem[12331] = 32'b11111011000111111101001100101000;
   assign mem[12332] = 32'b11111011000111101100111111101000;
   assign mem[12333] = 32'b00001000001111110111011000010000;
   assign mem[12334] = 32'b00001010100111010011000111010000;
   assign mem[12335] = 32'b11111110000101111100000001100110;
   assign mem[12336] = 32'b11111110010011110110100000000100;
   assign mem[12337] = 32'b00000010110110110100110001000000;
   assign mem[12338] = 32'b11111111101111011101010111000001;
   assign mem[12339] = 32'b11111111010011101111011111001000;
   assign mem[12340] = 32'b11110101100100010001110010100000;
   assign mem[12341] = 32'b00000000000000100100101001000101;
   assign mem[12342] = 32'b00000010000110111100111101101000;
   assign mem[12343] = 32'b11111100110011011001110101010000;
   assign mem[12344] = 32'b00000100011010110111001111110000;
   assign mem[12345] = 32'b11111010111001110100110111001000;
   assign mem[12346] = 32'b11111110100111011100101111101010;
   assign mem[12347] = 32'b00000100100001101101111010100000;
   assign mem[12348] = 32'b00000010110010100001111001010000;
   assign mem[12349] = 32'b11111001011100110001110011100000;
   assign mem[12350] = 32'b00001001011111110011001100010000;
   assign mem[12351] = 32'b00000000110100101011011111011111;
   assign mem[12352] = 32'b00000001000111101110010011111000;
   assign mem[12353] = 32'b11111110111011000111000000110010;
   assign mem[12354] = 32'b11111111010010100110010100010001;
   assign mem[12355] = 32'b11111000101001001010101100111000;
   assign mem[12356] = 32'b00000011011101111100101010111100;
   assign mem[12357] = 32'b11111111011100010110111101011101;
   assign mem[12358] = 32'b00000101101001000110111101111000;
   assign mem[12359] = 32'b11110101000100001001100110110000;
   assign mem[12360] = 32'b00000100011100010000101010010000;
   assign mem[12361] = 32'b11111100110111111101111101001100;
   assign mem[12362] = 32'b00000011000111000111001010011100;
   assign mem[12363] = 32'b11111001100111100010001111110000;
   assign mem[12364] = 32'b00000001011110001101100100011100;
   assign mem[12365] = 32'b11111101101101001001011010111100;
   assign mem[12366] = 32'b11110111010110011110000011100000;
   assign mem[12367] = 32'b00000101101000111010111111011000;
   assign mem[12368] = 32'b11111010001101000101110011110000;
   assign mem[12369] = 32'b11111101111110101000111101111000;
   assign mem[12370] = 32'b11111100100111011100000000101100;
   assign mem[12371] = 32'b00000010111000111010011011110000;
   assign mem[12372] = 32'b00000011011011111001110010001000;
   assign mem[12373] = 32'b00000011000001101111101111110100;
   assign mem[12374] = 32'b00000100010110101010111111011000;
   assign mem[12375] = 32'b11111101101100000111100110011100;
   assign mem[12376] = 32'b00000100110010110011110000110000;
   assign mem[12377] = 32'b11111010110101111110110110011000;
   assign mem[12378] = 32'b00000011101010011011010110111100;
   assign mem[12379] = 32'b11101001000000110001100111100000;
   assign mem[12380] = 32'b00000101000010010000000000001000;
   assign mem[12381] = 32'b11111110111001100110010100100000;
   assign mem[12382] = 32'b00000001010010000011011011000110;
   assign mem[12383] = 32'b00000010000101101000010011111000;
   assign mem[12384] = 32'b11110110001011001001010010000000;
   assign mem[12385] = 32'b11111101101101111110110101111000;
   assign mem[12386] = 32'b00000011110001100110100010011100;
   assign mem[12387] = 32'b00000011100011101011110001110000;
   assign mem[12388] = 32'b11111011111001010100010110011000;
   assign mem[12389] = 32'b11111111010111010011100011111010;
   assign mem[12390] = 32'b11111110100001000000001001110100;
   assign mem[12391] = 32'b11111100110001101011110101101100;
   assign mem[12392] = 32'b11111111110101000000110001111000;
   assign mem[12393] = 32'b11111111010010000010011010111011;
   assign mem[12394] = 32'b00000011111101101010101101000100;
   assign mem[12395] = 32'b00000010100011100001010110010100;
   assign mem[12396] = 32'b00000010000011100010011010110100;
   assign mem[12397] = 32'b11110111110101101100101001000000;
   assign mem[12398] = 32'b00000001000010111001101010111100;
   assign mem[12399] = 32'b00000101001000110110111000010000;
   assign mem[12400] = 32'b11111111101101000111001010111100;
   assign mem[12401] = 32'b11111011111110000101010110011000;
   assign mem[12402] = 32'b11111011010011100001100111111000;
   assign mem[12403] = 32'b00000000111001110101010011011010;
   assign mem[12404] = 32'b00000100010110110001110110001000;
   assign mem[12405] = 32'b00000100100110001000010010010000;
   assign mem[12406] = 32'b11111011101101101001100000111000;
   assign mem[12407] = 32'b11110100101110100101101010010000;
   assign mem[12408] = 32'b00000011111011100000001100100100;
   assign mem[12409] = 32'b00000011000001110101100001011100;
   assign mem[12410] = 32'b00000001001001000111101011001000;
   assign mem[12411] = 32'b11111011111001100011110101001000;
   assign mem[12412] = 32'b11111101101101101110111010111000;
   assign mem[12413] = 32'b00000000111010000010101000111110;
   assign mem[12414] = 32'b00000001101001101011000110000110;
   assign mem[12415] = 32'b00000000010000010011110010110111;
   assign mem[12416] = 32'b00000000010110010010101000000011;
   assign mem[12417] = 32'b11111111001111011100110011110110;
   assign mem[12418] = 32'b11111101011001110011001110001100;
   assign mem[12419] = 32'b11111111110101110110110001011011;
   assign mem[12420] = 32'b11111100101111000000010001011000;
   assign mem[12421] = 32'b00000000110011011101001010011011;
   assign mem[12422] = 32'b11111100101110111101101101100100;
   assign mem[12423] = 32'b11111101001000110000011001011100;
   assign mem[12424] = 32'b00000101010010000000101110000000;
   assign mem[12425] = 32'b11111110000111100010011111011000;
   assign mem[12426] = 32'b11111001000011000100101011011000;
   assign mem[12427] = 32'b00000010011011000100101011110100;
   assign mem[12428] = 32'b00000000101101001011100011100010;
   assign mem[12429] = 32'b11111111110010010011001010010101;
   assign mem[12430] = 32'b11111110101111010110100111011110;
   assign mem[12431] = 32'b11111100111010001100001110001000;
   assign mem[12432] = 32'b00000101101011100111111001011000;
   assign mem[12433] = 32'b11111101101011100101000110011000;
   assign mem[12434] = 32'b00000101010110111100110011010000;
   assign mem[12435] = 32'b11110000101011110010001010100000;
   assign mem[12436] = 32'b11110100010011111101000001100000;
   assign mem[12437] = 32'b00000011010101100000000111001000;
   assign mem[12438] = 32'b11111011111101000111100101001000;
   assign mem[12439] = 32'b00000001011011101010101111100110;
   assign mem[12440] = 32'b00000011100001001001010111010000;
   assign mem[12441] = 32'b00000101011111011111100111101000;
   assign mem[12442] = 32'b00001000001111001010100101100000;
   assign mem[12443] = 32'b11111100101110110010110011001100;
   assign mem[12444] = 32'b00000011001110111101110100111100;
   assign mem[12445] = 32'b11110101101011110101001101010000;
   assign mem[12446] = 32'b11111111110111011111000100011100;
   assign mem[12447] = 32'b00000000011110111100000111101101;
   assign mem[12448] = 32'b00000000111010010001010010111010;
   assign mem[12449] = 32'b11110101100100110010100000000000;
   assign mem[12450] = 32'b11111000101110001110010001100000;
   assign mem[12451] = 32'b11111110000011000110101100000000;
   assign mem[12452] = 32'b00000100110011011100010010001000;
   assign mem[12453] = 32'b00000010001011110110010111000100;
   assign mem[12454] = 32'b00000011011100100011100101110100;
   assign mem[12455] = 32'b00000100101011110000000001001000;
   assign mem[12456] = 32'b00000000110000000110110101101001;
   assign mem[12457] = 32'b11111010100101001100101010110000;
   assign mem[12458] = 32'b00000000100011110111101011110100;
   assign mem[12459] = 32'b11110111001101110001100010010000;
   assign mem[12460] = 32'b11111111000100001011001000110111;
   assign mem[12461] = 32'b11111010011100101001101010011000;
   assign mem[12462] = 32'b11111010101100010101011101011000;
   assign mem[12463] = 32'b00000101010100011001000101001000;
   assign mem[12464] = 32'b00000110101101010101101001000000;
   assign mem[12465] = 32'b11111101100011101111101110010000;
   assign mem[12466] = 32'b11111110101101100100000001110100;
   assign mem[12467] = 32'b11111010110010001011001101110000;
   assign mem[12468] = 32'b00000001101010101111100000110010;
   assign mem[12469] = 32'b00000010000001000100001110010100;
   assign mem[12470] = 32'b00000101111100000101010100100000;
   assign mem[12471] = 32'b11110101010010101011001001110000;
   assign mem[12472] = 32'b00001010101100101111011010110000;
   assign mem[12473] = 32'b11110010111011000000101100110000;
   assign mem[12474] = 32'b00000111010101001110000111010000;
   assign mem[12475] = 32'b11110101010111000011111001110000;
   assign mem[12476] = 32'b11111101100101011011011110000100;
   assign mem[12477] = 32'b00000110010110100100000111111000;
   assign mem[12478] = 32'b11111001111101110011101111010000;
   assign mem[12479] = 32'b11110110100010011110110000000000;
   assign mem[12480] = 32'b00000010111010111100100010110100;
   assign mem[12481] = 32'b00000010001100111110011011010100;
   assign mem[12482] = 32'b00000010111000101001110011011100;
   assign mem[12483] = 32'b11111111101110001000110101101010;
   assign mem[12484] = 32'b11111001000000100011000111011000;
   assign mem[12485] = 32'b11111110000100110001001000101010;
   assign mem[12486] = 32'b00000010101000101100000110000100;
   assign mem[12487] = 32'b00000110001110111010111011001000;
   assign mem[12488] = 32'b11111000000001101111011100011000;
   assign mem[12489] = 32'b00000100100111111100100101101000;
   assign mem[12490] = 32'b00001000110100100000001001110000;
   assign mem[12491] = 32'b11101111001100111111001010100000;
   assign mem[12492] = 32'b00001000101101010111110000110000;
   assign mem[12493] = 32'b11111110100111100100100011010010;
   assign mem[12494] = 32'b11111110011000110000011111101110;
   assign mem[12495] = 32'b11111111001101111100000111110010;
   assign mem[12496] = 32'b11111101100100100101100110110000;
   assign mem[12497] = 32'b00001100100011010101010010010000;
   assign mem[12498] = 32'b11110000001011011111110110100000;
   assign mem[12499] = 32'b00000000100001110101011001000100;
   assign mem[12500] = 32'b00000100011000110001010011000000;
   assign mem[12501] = 32'b11111111001000011100000001101111;
   assign mem[12502] = 32'b00000110101101010001001111100000;
   assign mem[12503] = 32'b11111000111101110000100001011000;
   assign mem[12504] = 32'b00000111101111010011101101111000;
   assign mem[12505] = 32'b11111001011001010110110001000000;
   assign mem[12506] = 32'b11111101110110001001100111100100;
   assign mem[12507] = 32'b00000111010111110101100011011000;
   assign mem[12508] = 32'b11111000011101100000101111001000;
   assign mem[12509] = 32'b11111011011111000110101111001000;
   assign mem[12510] = 32'b00000011001000010011110000111000;
   assign mem[12511] = 32'b11111010011100010110001011101000;
   assign mem[12512] = 32'b11111010101110110010100000001000;
   assign mem[12513] = 32'b00000010111111110001011011000000;
   assign mem[12514] = 32'b11111110011000001000110011011110;
   assign mem[12515] = 32'b00000001011000001101000100001100;
   assign mem[12516] = 32'b00000011000000010101111001011100;
   assign mem[12517] = 32'b00000110001010011101010101101000;
   assign mem[12518] = 32'b11111101100100011000000101110000;
   assign mem[12519] = 32'b00000001000101011010101001111000;
   assign mem[12520] = 32'b11110001000000000000011001010000;
   assign mem[12521] = 32'b00000010010000001011111000001000;
   assign mem[12522] = 32'b00000001111111010010011000010100;
   assign mem[12523] = 32'b00000001100001010101011101000010;
   assign mem[12524] = 32'b11111001101011111000110010110000;
   assign mem[12525] = 32'b00000000001111101010001010010011;
   assign mem[12526] = 32'b00000111000010100010000101011000;
   assign mem[12527] = 32'b00000100011100111010111010110000;
   assign mem[12528] = 32'b00001000001101110010110100000000;
   assign mem[12529] = 32'b11101110100101100111100111000000;
   assign mem[12530] = 32'b11110001010101111100010101100000;
   assign mem[12531] = 32'b00000010011101000111111100100000;
   assign mem[12532] = 32'b11111111001011100100010111100110;
   assign mem[12533] = 32'b00000100010010110111010001110000;
   assign mem[12534] = 32'b00000101011111100101110101010000;
   assign mem[12535] = 32'b00000001100110110111010001010100;
   assign mem[12536] = 32'b11111100101001111110000110100100;
   assign mem[12537] = 32'b00001001000111000011101011000000;
   assign mem[12538] = 32'b00000100101110111000100001101000;
   assign mem[12539] = 32'b11111001110111010011001011100000;
   assign mem[12540] = 32'b00000011010001100111111101010100;
   assign mem[12541] = 32'b11111110001100001000000111011110;
   assign mem[12542] = 32'b00000011001001101100011111101000;
   assign mem[12543] = 32'b11111100000110010100101111101000;
   assign mem[12544] = 32'b00000100100100100001011011100000;
   assign mem[12545] = 32'b11111001011001000011111010101000;
   assign mem[12546] = 32'b00000100011111111111000101111000;
   assign mem[12547] = 32'b00000011101100111001111011001100;
   assign mem[12548] = 32'b11110001011000111001110001010000;
   assign mem[12549] = 32'b11111101010110100111001110011000;
   assign mem[12550] = 32'b11111111111101110110010011011100;
   assign mem[12551] = 32'b11111010001000110101010111011000;
   assign mem[12552] = 32'b00001100010000010011111101000000;
   assign mem[12553] = 32'b11101101010101011100111000100000;
   assign mem[12554] = 32'b11111001111011110101110100100000;
   assign mem[12555] = 32'b00000010100101001010100011011100;
   assign mem[12556] = 32'b11101100111001000100011000000000;
   assign mem[12557] = 32'b11111110100010010000100100111110;
   assign mem[12558] = 32'b00000110001010101000111110101000;
   assign mem[12559] = 32'b11111000100110010100101100101000;
   assign mem[12560] = 32'b00000101010110100010111010101000;
   assign mem[12561] = 32'b11110101000000111000110100100000;
   assign mem[12562] = 32'b00001101000001100110101111010000;
   assign mem[12563] = 32'b11111000110111111111011000110000;
   assign mem[12564] = 32'b11111110010000100101010010110110;
   assign mem[12565] = 32'b00000000011111101001111101010100;
   assign mem[12566] = 32'b00000010110001000101001101011000;
   assign mem[12567] = 32'b11111111101000111000111011111101;
   assign mem[12568] = 32'b11111011101000011011100100110000;
   assign mem[12569] = 32'b00000001101111011100011000011110;
   assign mem[12570] = 32'b00001000101110101010110001010000;
   assign mem[12571] = 32'b11110010110001001011101101110000;
   assign mem[12572] = 32'b11111111000101001111100011000011;
   assign mem[12573] = 32'b11110110110101001111111000100000;
   assign mem[12574] = 32'b00000100110011001100001010111000;
   assign mem[12575] = 32'b11101010000111010011010011100000;
   assign mem[12576] = 32'b00000100000100110011111110111000;
   assign mem[12577] = 32'b00001000101111000010001110010000;
   assign mem[12578] = 32'b11111101100100000001101000000000;
   assign mem[12579] = 32'b00000001001011010001010011111100;
   assign mem[12580] = 32'b11111101000111000000010100001100;
   assign mem[12581] = 32'b00000000011010011010001101111010;
   assign mem[12582] = 32'b00010001000010011010010011000000;
   assign mem[12583] = 32'b11101000000101011100101001100000;
   assign mem[12584] = 32'b11111100011001100010111000010100;
   assign mem[12585] = 32'b00000100110000110010011100101000;
   assign mem[12586] = 32'b11110001110101101110101010100000;
   assign mem[12587] = 32'b00000101011111000100011111011000;
   assign mem[12588] = 32'b11111100100010011101100000110100;
   assign mem[12589] = 32'b11111101000010100100010010111000;
   assign mem[12590] = 32'b00000001100000110001110010110100;
   assign mem[12591] = 32'b00000001010100101111011011111010;
   assign mem[12592] = 32'b11111011100101101100111011000000;
   assign mem[12593] = 32'b00000100001001001100111111101000;
   assign mem[12594] = 32'b11111101000000001010101011010000;
   assign mem[12595] = 32'b00000100101100101011011001000000;
   assign mem[12596] = 32'b00000101110000110101100110100000;
   assign mem[12597] = 32'b11111011110001101100110110100000;
   assign mem[12598] = 32'b00000100010001101000000010110000;
   assign mem[12599] = 32'b00000000001100110111100111110100;
   assign mem[12600] = 32'b11111011111001010011011001010000;
   assign mem[12601] = 32'b00000000010001111010010101000111;
   assign mem[12602] = 32'b00000101111000010111101100110000;
   assign mem[12603] = 32'b00000010100100010101001101011000;
   assign mem[12604] = 32'b00000001001111011110000111010110;
   assign mem[12605] = 32'b00000001010010100011010110000100;
   assign mem[12606] = 32'b00000000000011010111011000110111;
   assign mem[12607] = 32'b00000011110001101000011100110100;
   assign mem[12608] = 32'b11101100101100000011001010100000;
   assign mem[12609] = 32'b00000001100000100100110110011110;
   assign mem[12610] = 32'b11111001110001110011000010100000;
   assign mem[12611] = 32'b11111100101101100000001100111000;
   assign mem[12612] = 32'b11111000100100110111011110010000;
   assign mem[12613] = 32'b00000110111010110101100011101000;
   assign mem[12614] = 32'b11110101000101000001111110110000;
   assign mem[12615] = 32'b00001000010101111100001111110000;
   assign mem[12616] = 32'b00000100011001011110001101000000;
   assign mem[12617] = 32'b11111101110001100011000111000100;
   assign mem[12618] = 32'b00000110000111100101101001100000;
   assign mem[12619] = 32'b11111010011110111000111000101000;
   assign mem[12620] = 32'b00000011111101110110111110000000;
   assign mem[12621] = 32'b11111100100001100101111000011000;
   assign mem[12622] = 32'b00000110000100110000100000111000;
   assign mem[12623] = 32'b11111101100111010010001001011000;
   assign mem[12624] = 32'b11111010011111000010111001000000;
   assign mem[12625] = 32'b00000011011110000011111011010000;
   assign mem[12626] = 32'b11111001001011111110100011010000;
   assign mem[12627] = 32'b11111011111100010110111101100000;
   assign mem[12628] = 32'b00000010001000101000011111011000;
   assign mem[12629] = 32'b11110100110100101001101100010000;
   assign mem[12630] = 32'b00000001001111010001011010010000;
   assign mem[12631] = 32'b11111110010010110010000010110100;
   assign mem[12632] = 32'b00000001011110110100001100001110;
   assign mem[12633] = 32'b00000001011101001111111110001010;
   assign mem[12634] = 32'b11111111100111001001000111101111;
   assign mem[12635] = 32'b00000000000111110010111110000100;
   assign mem[12636] = 32'b00000001011100111110010000001100;
   assign mem[12637] = 32'b11111111011010111001011011000101;
   assign mem[12638] = 32'b11111101011110100101010111111000;
   assign mem[12639] = 32'b00000000001110110001110100101001;
   assign mem[12640] = 32'b00000001100011011011110111000010;
   assign mem[12641] = 32'b11111101011111111000000001101100;
   assign mem[12642] = 32'b11111111000111110100101010011010;
   assign mem[12643] = 32'b11111110000011111001000000101100;
   assign mem[12644] = 32'b00000101100110101100111110001000;
   assign mem[12645] = 32'b11111101110110010000100100101000;
   assign mem[12646] = 32'b00000011001011101110111010010000;
   assign mem[12647] = 32'b00000001111111000110010100111100;
   assign mem[12648] = 32'b11110001111101101001011110010000;
   assign mem[12649] = 32'b00000011000000101000111011100100;
   assign mem[12650] = 32'b11111001000111011011001000101000;
   assign mem[12651] = 32'b11111101110010110110000110110000;
   assign mem[12652] = 32'b00001110011000011010110001000000;
   assign mem[12653] = 32'b11111100101100100010111111100100;
   assign mem[12654] = 32'b11111100110101010011000001110100;
   assign mem[12655] = 32'b11111010100000110000011010101000;
   assign mem[12656] = 32'b00000000000100100110010100001011;
   assign mem[12657] = 32'b00001001001110101000100011000000;
   assign mem[12658] = 32'b11110100100001110110000101000000;
   assign mem[12659] = 32'b11111110010000101100010010111000;
   assign mem[12660] = 32'b00000011010110101001000001111000;
   assign mem[12661] = 32'b00000000000001100101111011111101;
   assign mem[12662] = 32'b11111101011001000101011001011000;
   assign mem[12663] = 32'b00000011001010101001010101000100;
   assign mem[12664] = 32'b11111111111001101111110110111101;
   assign mem[12665] = 32'b00000000001110111010001011110100;
   assign mem[12666] = 32'b00000010101010100111010010111000;
   assign mem[12667] = 32'b00000001100100001011100011001100;
   assign mem[12668] = 32'b00000011000000111000010111001000;
   assign mem[12669] = 32'b11111100110010100110000011100100;
   assign mem[12670] = 32'b00000001011101010000000101010100;
   assign mem[12671] = 32'b00001011111111011001010000110000;
   assign mem[12672] = 32'b11101110110011111100111100000000;
   assign mem[12673] = 32'b11111110110001101111111001100010;
   assign mem[12674] = 32'b11110111100001101000110110000000;
   assign mem[12675] = 32'b00000001010100010000010110001010;
   assign mem[12676] = 32'b11111100010011111011100010010100;
   assign mem[12677] = 32'b11111000010110000110011010101000;
   assign mem[12678] = 32'b00001011010001010110111100110000;
   assign mem[12679] = 32'b11111100110111000001100110001000;
   assign mem[12680] = 32'b00001001101010001001101101110000;
   assign mem[12681] = 32'b11111101001010000000001110000100;
   assign mem[12682] = 32'b00000111110100000010101111101000;
   assign mem[12683] = 32'b11110111001100110111010010000000;
   assign mem[12684] = 32'b00000011111000011010101101101100;
   assign mem[12685] = 32'b11111001111111011101011100111000;
   assign mem[12686] = 32'b00000001101001000111101111110010;
   assign mem[12687] = 32'b00000111011100000101000100011000;
   assign mem[12688] = 32'b11111101111011011110011100001000;
   assign mem[12689] = 32'b11101101110011100100110000000000;
   assign mem[12690] = 32'b11111011000010110111011101101000;
   assign mem[12691] = 32'b00000010101111100101000011100100;
   assign mem[12692] = 32'b00000001110000000100101010000010;
   assign mem[12693] = 32'b11111011101110010010000000011000;
   assign mem[12694] = 32'b00000100010011111001101001000000;
   assign mem[12695] = 32'b00000001111011011000110010001000;
   assign mem[12696] = 32'b11111101110100010010101000010000;
   assign mem[12697] = 32'b00000001011011100001010110001000;
   assign mem[12698] = 32'b00000000100100001110101101100101;
   assign mem[12699] = 32'b11101011111111111111100010000000;
   assign mem[12700] = 32'b00000111110010011101011011110000;
   assign mem[12701] = 32'b11111101000110001100100110110100;
   assign mem[12702] = 32'b00000100010100111101101101100000;
   assign mem[12703] = 32'b11111111000000111101010010011111;
   assign mem[12704] = 32'b00000010000010010011101011010000;
   assign mem[12705] = 32'b11111000100100101101001110100000;
   assign mem[12706] = 32'b00000010111011110000100000110100;
   assign mem[12707] = 32'b00000111001011000100110010111000;
   assign mem[12708] = 32'b11111000101100100000001001110000;
   assign mem[12709] = 32'b11111000001000101011010111011000;
   assign mem[12710] = 32'b11111110101001111000101011111100;
   assign mem[12711] = 32'b11101110110001001001001111000000;
   assign mem[12712] = 32'b11111110101010111110100110000000;
   assign mem[12713] = 32'b00000011100000001110100100001000;
   assign mem[12714] = 32'b11110110111011011110101110110000;
   assign mem[12715] = 32'b11111110000001101010011011010000;
   assign mem[12716] = 32'b00000010010110000101111001010000;
   assign mem[12717] = 32'b00000100011100010100101110111000;
   assign mem[12718] = 32'b11111111111110100010110111100011;
   assign mem[12719] = 32'b11111101001101101111101001010000;
   assign mem[12720] = 32'b11111110110101100101000000010000;
   assign mem[12721] = 32'b11111000100101001110001111100000;
   assign mem[12722] = 32'b11111000001011110001100100101000;
   assign mem[12723] = 32'b00000000110001000000101100011100;
   assign mem[12724] = 32'b11111101100100100010011110101100;
   assign mem[12725] = 32'b00000010010100110101101001011100;
   assign mem[12726] = 32'b00000010000001111010101101111000;
   assign mem[12727] = 32'b11111101110111000100011011010000;
   assign mem[12728] = 32'b00000001100000100010011010100000;
   assign mem[12729] = 32'b00000001001000110000010000000110;
   assign mem[12730] = 32'b00000010000111000000111000101100;
   assign mem[12731] = 32'b11111110001111110100110111010010;
   assign mem[12732] = 32'b00000100110111001110010010010000;
   assign mem[12733] = 32'b00000001111110000011010100011100;
   assign mem[12734] = 32'b11111101010101110011010101100100;
   assign mem[12735] = 32'b00000010111111100001010001011000;
   assign mem[12736] = 32'b11111110011011111001000011011010;
   assign mem[12737] = 32'b11111011010000010000010111010000;
   assign mem[12738] = 32'b00000001010010111010011010011000;
   assign mem[12739] = 32'b11110000001011100001010000110000;
   assign mem[12740] = 32'b11110010110011000110000101010000;
   assign mem[12741] = 32'b00000000000111111101101000110010;
   assign mem[12742] = 32'b00000001111100000111101101111010;
   assign mem[12743] = 32'b00001000110001100100001100110000;
   assign mem[12744] = 32'b11101111010011010000010111100000;
   assign mem[12745] = 32'b00000001001100010110100110111100;
   assign mem[12746] = 32'b00000010000101001011010111001100;
   assign mem[12747] = 32'b11111000000001110010001111011000;
   assign mem[12748] = 32'b00000010110100000000111110011000;
   assign mem[12749] = 32'b11111000101011010001100101000000;
   assign mem[12750] = 32'b11111001001111110101000100001000;
   assign mem[12751] = 32'b11111110000011010001101101001110;
   assign mem[12752] = 32'b11111011101100011001011100001000;
   assign mem[12753] = 32'b00000011101101101010101000101100;
   assign mem[12754] = 32'b11111000101011100110010110011000;
   assign mem[12755] = 32'b00000001110010010100100100100010;
   assign mem[12756] = 32'b00000110000111111011110101111000;
   assign mem[12757] = 32'b11110111011001110000110010100000;
   assign mem[12758] = 32'b00000101111101100000000111111000;
   assign mem[12759] = 32'b11111000010111101000001101011000;
   assign mem[12760] = 32'b11110111010111000010111000110000;
   assign mem[12761] = 32'b00000000100111111101100001101110;
   assign mem[12762] = 32'b00010011110111110010110010100000;
   assign mem[12763] = 32'b11110010110001000011111000010000;
   assign mem[12764] = 32'b00000011001010000111110011001000;
   assign mem[12765] = 32'b00000010110110101001100001110100;
   assign mem[12766] = 32'b11111011110001111100010111001000;
   assign mem[12767] = 32'b00001001011110010000010000010000;
   assign mem[12768] = 32'b11110100110000010001110110010000;
   assign mem[12769] = 32'b11111010011011110110110111101000;
   assign mem[12770] = 32'b00000000101100011000001000111011;
   assign mem[12771] = 32'b11111101100000110110010010010100;
   assign mem[12772] = 32'b00010011010011010100001101000000;
   assign mem[12773] = 32'b11111101110100100101001111100100;
   assign mem[12774] = 32'b00001010000010000111110101000000;
   assign mem[12775] = 32'b11111111011111101010111011000111;
   assign mem[12776] = 32'b00000001000101000111101001001000;
   assign mem[12777] = 32'b00001111111110100010111100010000;
   assign mem[12778] = 32'b11110000010010000100100000010000;
   assign mem[12779] = 32'b11111001010000100100101111110000;
   assign mem[12780] = 32'b00000001101100101100000101000100;
   assign mem[12781] = 32'b11111011111010010100110010010000;
   assign mem[12782] = 32'b00000101101011100001011111010000;
   assign mem[12783] = 32'b11110111111100010100000110000000;
   assign mem[12784] = 32'b00000100001111100010001000010000;
   assign mem[12785] = 32'b11111110100011110010110011000100;
   assign mem[12786] = 32'b11111101000011000001110100010000;
   assign mem[12787] = 32'b00000000101011001011010001011010;
   assign mem[12788] = 32'b11110010000000101001001110110000;
   assign mem[12789] = 32'b00000110011011111101111101010000;
   assign mem[12790] = 32'b00001000111011000100011101100000;
   assign mem[12791] = 32'b11110001010010000011011001110000;
   assign mem[12792] = 32'b11110111001011110111000101010000;
   assign mem[12793] = 32'b11111101111100010100000111111000;
   assign mem[12794] = 32'b11111111101110001001010110110011;
   assign mem[12795] = 32'b11111110100000101001011100100110;
   assign mem[12796] = 32'b11111101000101100011000100110100;
   assign mem[12797] = 32'b00000110100111110100010111011000;
   assign mem[12798] = 32'b11111011110000000010111100101000;
   assign mem[12799] = 32'b11111010101101011101101111000000;
   assign mem[12800] = 32'b00000000001001001001110101010101;
   assign mem[12801] = 32'b11111010011110101001110101110000;
   assign mem[12802] = 32'b00000010000001001001111110000100;
   assign mem[12803] = 32'b00000001101110110001001101100110;
   assign mem[12804] = 32'b11111101000001111010000111110000;
   assign mem[12805] = 32'b11111111011011110100111000110110;
   assign mem[12806] = 32'b00000010001100000010100010101100;
   assign mem[12807] = 32'b11111111001000011011000000000101;
   assign mem[12808] = 32'b11111100011011000000110111111000;
   assign mem[12809] = 32'b00000000100010111100001011100000;
   assign mem[12810] = 32'b11111000010111011001000001011000;
   assign mem[12811] = 32'b11111110000101111111111111010110;
   assign mem[12812] = 32'b11111101001110010101111100100100;
   assign mem[12813] = 32'b11111100010000011001011111101100;
   assign mem[12814] = 32'b00000001010111001110111001001010;
   assign mem[12815] = 32'b00000000010011101010100001010110;
   assign mem[12816] = 32'b11111111011111111111110100010110;
   assign mem[12817] = 32'b00001001001100100000100001100000;
   assign mem[12818] = 32'b11111110001001010001000111100000;
   assign mem[12819] = 32'b00000000011000100000100000000001;
   assign mem[12820] = 32'b00000110000011000111011111011000;
   assign mem[12821] = 32'b11110110111011101111010000100000;
   assign mem[12822] = 32'b11111001101000110001100001110000;
   assign mem[12823] = 32'b00000001001001011010100111000010;
   assign mem[12824] = 32'b00000001001011011010100010101110;
   assign mem[12825] = 32'b11111110110100111000001010111010;
   assign mem[12826] = 32'b00000010011010111011010011011000;
   assign mem[12827] = 32'b11110010010010011101011001010000;
   assign mem[12828] = 32'b00001010010101000011011101010000;
   assign mem[12829] = 32'b00000010100001001001000110000100;
   assign mem[12830] = 32'b11111101100001000100110111101100;
   assign mem[12831] = 32'b00001010001110010111100001110000;
   assign mem[12832] = 32'b11111101000011000011001110111000;
   assign mem[12833] = 32'b11111111010000101101010111110111;
   assign mem[12834] = 32'b00000001101011000110010000111010;
   assign mem[12835] = 32'b11111111110001110110110111101010;
   assign mem[12836] = 32'b00000010000011010100110000000000;
   assign mem[12837] = 32'b11111100011111011000100100001000;
   assign mem[12838] = 32'b11111111000011111001111010001000;
   assign mem[12839] = 32'b11111100101010111011000011111000;
   assign mem[12840] = 32'b00000001011001011100011001110110;
   assign mem[12841] = 32'b00000111111011011111000010100000;
   assign mem[12842] = 32'b11111101011000111110101000010100;
   assign mem[12843] = 32'b11111110001001110110011011010010;
   assign mem[12844] = 32'b00000110100001010110011101111000;
   assign mem[12845] = 32'b00000011010111011000110100010100;
   assign mem[12846] = 32'b11111111111100010111011110110001;
   assign mem[12847] = 32'b00000100111100101101001001001000;
   assign mem[12848] = 32'b11110101101110111110001000000000;
   assign mem[12849] = 32'b11111111111001100100011010111000;
   assign mem[12850] = 32'b00010000000011010100101010100000;
   assign mem[12851] = 32'b11111101001100111111000000101100;
   assign mem[12852] = 32'b00000111111101000011011011010000;
   assign mem[12853] = 32'b00000001011010000111011110010000;
   assign mem[12854] = 32'b11110001101111001001010011110000;
   assign mem[12855] = 32'b11111000000000101110010100101000;
   assign mem[12856] = 32'b11111001101011001001110011110000;
   assign mem[12857] = 32'b11111100011110100100001000100100;
   assign mem[12858] = 32'b00000100011001011100000101011000;
   assign mem[12859] = 32'b11110010001110100110110001000000;
   assign mem[12860] = 32'b00000100010101010101101011111000;
   assign mem[12861] = 32'b00001011101000100011101011110000;
   assign mem[12862] = 32'b00000010111000010110100111101000;
   assign mem[12863] = 32'b11111010100001010101011101100000;
   assign mem[12864] = 32'b00000001001010000001010101011100;
   assign mem[12865] = 32'b11110101001100010010000001010000;
   assign mem[12866] = 32'b11111101100010011011000010011100;
   assign mem[12867] = 32'b11111111111001010111101011101111;
   assign mem[12868] = 32'b00000010100010010001010010011100;
   assign mem[12869] = 32'b11111101100000001010010011101000;
   assign mem[12870] = 32'b11110110100101111001101111000000;
   assign mem[12871] = 32'b00001001101011101110001110100000;
   assign mem[12872] = 32'b00000011000010010100101101101000;
   assign mem[12873] = 32'b11110000101010010101111010110000;
   assign mem[12874] = 32'b00000100101001011110011111010000;
   assign mem[12875] = 32'b00000001011010000011100001111110;
   assign mem[12876] = 32'b11111110101010110011100101011010;
   assign mem[12877] = 32'b11111100111010111101111001110100;
   assign mem[12878] = 32'b00000011110011101000110111101000;
   assign mem[12879] = 32'b11111101100001110111111000010100;
   assign mem[12880] = 32'b11110100110100011100110001110000;
   assign mem[12881] = 32'b00001001111110001100111010000000;
   assign mem[12882] = 32'b11101011101110011011110010100000;
   assign mem[12883] = 32'b00001001000110100011010001110000;
   assign mem[12884] = 32'b00000001011100010000101000100100;
   assign mem[12885] = 32'b00000100111101011000000100001000;
   assign mem[12886] = 32'b11111011101101111011111110011000;
   assign mem[12887] = 32'b00000011011110111100010000011100;
   assign mem[12888] = 32'b11110111010000111010000000010000;
   assign mem[12889] = 32'b11111111011010101100110010010110;
   assign mem[12890] = 32'b00000101101011101000000000010000;
   assign mem[12891] = 32'b00000110100101110110111000000000;
   assign mem[12892] = 32'b00000110101000001001001001010000;
   assign mem[12893] = 32'b11111100100011110100110001000000;
   assign mem[12894] = 32'b00000000001010011111010101010100;
   assign mem[12895] = 32'b11111010010010110001010100011000;
   assign mem[12896] = 32'b00000001000111100000001001110110;
   assign mem[12897] = 32'b11111111101001110100000010000011;
   assign mem[12898] = 32'b11111110001011001110000110101110;
   assign mem[12899] = 32'b11111101000110010001010000001100;
   assign mem[12900] = 32'b11111111100011010011001010110100;
   assign mem[12901] = 32'b00001111001101100000001110010000;
   assign mem[12902] = 32'b11111111100000001000100110011111;
   assign mem[12903] = 32'b00000001010011101111100001011100;
   assign mem[12904] = 32'b11111001010110110100100010010000;
   assign mem[12905] = 32'b00000101010100100110110011000000;
   assign mem[12906] = 32'b11111011101100111011111000110000;
   assign mem[12907] = 32'b11111101111010100110001110101100;
   assign mem[12908] = 32'b00000000001110010000010111111000;
   assign mem[12909] = 32'b11111010100011001111101100101000;
   assign mem[12910] = 32'b00000000101001001111111010101100;
   assign mem[12911] = 32'b00000001000011110010011110110100;
   assign mem[12912] = 32'b11111011001101000111101110010000;
   assign mem[12913] = 32'b00000101011101010101101100111000;
   assign mem[12914] = 32'b11111111001011001110011001000100;
   assign mem[12915] = 32'b00000010111010010000101000110100;
   assign mem[12916] = 32'b00000000111110010110000011100101;
   assign mem[12917] = 32'b11111000010000000000001101011000;
   assign mem[12918] = 32'b11111101011001110110010111100100;
   assign mem[12919] = 32'b11111111011011100001001111000000;
   assign mem[12920] = 32'b11111100110101111101110001110100;
   assign mem[12921] = 32'b00000001110011011000001010100100;
   assign mem[12922] = 32'b11110110001011111010011111010000;
   assign mem[12923] = 32'b00010010101011100100101100100000;
   assign mem[12924] = 32'b11110010111000001011011011010000;
   assign mem[12925] = 32'b00000111101111011100101001111000;
   assign mem[12926] = 32'b11110100111010111010001110110000;
   assign mem[12927] = 32'b11110100101001100000000010100000;
   assign mem[12928] = 32'b11111101011011111101000111011000;
   assign mem[12929] = 32'b00000010101101000011001111011000;
   assign mem[12930] = 32'b11110110000101010010011010000000;
   assign mem[12931] = 32'b00000110100010111100111011011000;
   assign mem[12932] = 32'b11100110011110010000101100000000;
   assign mem[12933] = 32'b00010100110000001000001110100000;
   assign mem[12934] = 32'b11111001111100101000100110100000;
   assign mem[12935] = 32'b00000111111000011101110011000000;
   assign mem[12936] = 32'b11111001111000100000000111110000;
   assign mem[12937] = 32'b11111011100011001000111000110000;
   assign mem[12938] = 32'b11101011001100110011111000100000;
   assign mem[12939] = 32'b00000010101001100001011111111100;
   assign mem[12940] = 32'b00000011001001110011101101010000;
   assign mem[12941] = 32'b00000100111111100001000011100000;
   assign mem[12942] = 32'b00000100100000101101110101110000;
   assign mem[12943] = 32'b00000001010100110010110101000100;
   assign mem[12944] = 32'b00000000001111111000011011000000;
   assign mem[12945] = 32'b00000010010100011100110110110100;
   assign mem[12946] = 32'b00000010010011011001110000110000;
   assign mem[12947] = 32'b11111100100110111110010111110000;
   assign mem[12948] = 32'b11111001111010010000000000000000;
   assign mem[12949] = 32'b00000101110011011111100100011000;
   assign mem[12950] = 32'b00000100111000101110011011011000;
   assign mem[12951] = 32'b11111111001101011111110111011000;
   assign mem[12952] = 32'b00000011011000111001000110101000;
   assign mem[12953] = 32'b11111000111101100110011011001000;
   assign mem[12954] = 32'b11110100110010000001100001110000;
   assign mem[12955] = 32'b11111000101111101100000011011000;
   assign mem[12956] = 32'b11111110011111111010000000001010;
   assign mem[12957] = 32'b00000100100001100101000111111000;
   assign mem[12958] = 32'b11111110010001000011000110001000;
   assign mem[12959] = 32'b11111101110010011111101010101100;
   assign mem[12960] = 32'b00000001011101000000110111110010;
   assign mem[12961] = 32'b00000011011101100010111001011100;
   assign mem[12962] = 32'b00000011000000111000101101101000;
   assign mem[12963] = 32'b11111110000101111111001001111100;
   assign mem[12964] = 32'b00000011100101111110000000100100;
   assign mem[12965] = 32'b11111111111001111000010101100010;
   assign mem[12966] = 32'b11111100110110101100110100101100;
   assign mem[12967] = 32'b11111101000001010111010111010100;
   assign mem[12968] = 32'b11111111000101110000101101110110;
   assign mem[12969] = 32'b11111101101110001001100101000100;
   assign mem[12970] = 32'b00000101001000100100100001110000;
   assign mem[12971] = 32'b11110011101000010110101110110000;
   assign mem[12972] = 32'b00000001010101001000100101011110;
   assign mem[12973] = 32'b00000011101101010000000110100000;
   assign mem[12974] = 32'b11110101110110011010111010110000;
   assign mem[12975] = 32'b11111111100010111010110101111000;
   assign mem[12976] = 32'b00000000111011001000010101011100;
   assign mem[12977] = 32'b11111011010011001000100101010000;
   assign mem[12978] = 32'b00000100000101011100100100101000;
   assign mem[12979] = 32'b11111000110010010111111101100000;
   assign mem[12980] = 32'b00000001000001110111101100101010;
   assign mem[12981] = 32'b00000110111110101101111110100000;
   assign mem[12982] = 32'b11111010111001110111010111001000;
   assign mem[12983] = 32'b11111111001111110000001000100000;
   assign mem[12984] = 32'b00000111101110000111010101110000;
   assign mem[12985] = 32'b11111011000001101100000001101000;
   assign mem[12986] = 32'b00000011111001100111011111111100;
   assign mem[12987] = 32'b00000010110000110110011100101100;
   assign mem[12988] = 32'b11110011001100011110111010000000;
   assign mem[12989] = 32'b00000010001100011110001100000100;
   assign mem[12990] = 32'b11111011101110001111101010001000;
   assign mem[12991] = 32'b00000110010111010011101101010000;
   assign mem[12992] = 32'b11111110110110001011011000110000;
   assign mem[12993] = 32'b11111001110110011101000110101000;
   assign mem[12994] = 32'b00000111100100010110000010000000;
   assign mem[12995] = 32'b00000100101011101110001111001000;
   assign mem[12996] = 32'b11110011101000110000111100000000;
   assign mem[12997] = 32'b00001000100001010111001011010000;
   assign mem[12998] = 32'b11110100001001101000111000000000;
   assign mem[12999] = 32'b11111101011101110011001101000000;
   assign mem[13000] = 32'b00000111111101110101101101111000;
   assign mem[13001] = 32'b00000001101110011110110010100000;
   assign mem[13002] = 32'b00000000110010111100011001000101;
   assign mem[13003] = 32'b11111110111101100010111101011010;
   assign mem[13004] = 32'b11110100001010001011101101000000;
   assign mem[13005] = 32'b11111000111111111011101100000000;
   assign mem[13006] = 32'b00000100100110000000011001100000;
   assign mem[13007] = 32'b11111110101110011101101001101110;
   assign mem[13008] = 32'b00000001010100000100110010001110;
   assign mem[13009] = 32'b11111001001001001011011011010000;
   assign mem[13010] = 32'b11111101000110001010110010011000;
   assign mem[13011] = 32'b00001011101100001000100001010000;
   assign mem[13012] = 32'b11110000111100101111111000010000;
   assign mem[13013] = 32'b00000001101010000010100111011010;
   assign mem[13014] = 32'b11111100010010001010001100011100;
   assign mem[13015] = 32'b00000101000111100001101111010000;
   assign mem[13016] = 32'b11110001100101101101111111100000;
   assign mem[13017] = 32'b00000000010101100010111001100111;
   assign mem[13018] = 32'b11111101101010100011011001000000;
   assign mem[13019] = 32'b11111101000011010111011000000100;
   assign mem[13020] = 32'b00000001010010110011110010100110;
   assign mem[13021] = 32'b00000000111100000011100111010011;
   assign mem[13022] = 32'b00001000100110100001111001010000;
   assign mem[13023] = 32'b11111101001100100011010011101000;
   assign mem[13024] = 32'b00000001100100001011011101010100;
   assign mem[13025] = 32'b11111111110001101111010100001010;
   assign mem[13026] = 32'b00000000001000011011111101110000;
   assign mem[13027] = 32'b11111011011110011100110001011000;
   assign mem[13028] = 32'b11111011001100011011011000100000;
   assign mem[13029] = 32'b00000001101000010011000100000100;
   assign mem[13030] = 32'b00000100010111101101101110100000;
   assign mem[13031] = 32'b11101111110111000000001110000000;
   assign mem[13032] = 32'b00001010110001111011001111010000;
   assign mem[13033] = 32'b00000001001000110010101001011110;
   assign mem[13034] = 32'b11111011001001000001010100010000;
   assign mem[13035] = 32'b11111101101000011101101001111000;
   assign mem[13036] = 32'b11111011011011100011000000101000;
   assign mem[13037] = 32'b11110100010101110001101110110000;
   assign mem[13038] = 32'b00000101010010100110000111001000;
   assign mem[13039] = 32'b11111101011001010110101101000000;
   assign mem[13040] = 32'b00000001101000100001001010010000;
   assign mem[13041] = 32'b11110111111110101001001100000000;
   assign mem[13042] = 32'b00000001010110011101111111111000;
   assign mem[13043] = 32'b00000101001001001000010000001000;
   assign mem[13044] = 32'b11110011010001000010101111000000;
   assign mem[13045] = 32'b00000000010000101111000100010111;
   assign mem[13046] = 32'b11111110000101100001101010100110;
   assign mem[13047] = 32'b11101101000110100111001011100000;
   assign mem[13048] = 32'b00000101110100100110110111011000;
   assign mem[13049] = 32'b11111110100010001001011010111110;
   assign mem[13050] = 32'b11111110011011100000001001111000;
   assign mem[13051] = 32'b11111100111101110100111011100100;
   assign mem[13052] = 32'b00001100100011011110011111000000;
   assign mem[13053] = 32'b11101100000001010010110001100000;
   assign mem[13054] = 32'b00000111110001010000101101101000;
   assign mem[13055] = 32'b00000100001000000101000000101000;
   assign mem[13056] = 32'b11111100100001111101111000001000;
   assign mem[13057] = 32'b11111100101101000110010101110000;
   assign mem[13058] = 32'b11111001101000100010000110001000;
   assign mem[13059] = 32'b11111010010000001010100010100000;
   assign mem[13060] = 32'b00000010111110001100100001010100;
   assign mem[13061] = 32'b11111011001111011111110011000000;
   assign mem[13062] = 32'b00001100101111110010110011100000;
   assign mem[13063] = 32'b00000001011000010100001101111110;
   assign mem[13064] = 32'b11111001110000100000010101011000;
   assign mem[13065] = 32'b11110100100011010101101111010000;
   assign mem[13066] = 32'b00000000000001101111100011111011;
   assign mem[13067] = 32'b11101010001001100111101100000000;
   assign mem[13068] = 32'b11111101011000101001000010111100;
   assign mem[13069] = 32'b11110001000011101001110110110000;
   assign mem[13070] = 32'b11101101101111001010001100000000;
   assign mem[13071] = 32'b00000110010111000011111111111000;
   assign mem[13072] = 32'b11111111001111100011110101011000;
   assign mem[13073] = 32'b00000010010110111001011101001000;
   assign mem[13074] = 32'b00000011000001101000011110110000;
   assign mem[13075] = 32'b00000110111010110010001110000000;
   assign mem[13076] = 32'b11101110010010111101100010000000;
   assign mem[13077] = 32'b00000011101111101110011000000000;
   assign mem[13078] = 32'b00000001110101011110100000101100;
   assign mem[13079] = 32'b00000100101100111100010010101000;
   assign mem[13080] = 32'b00000011101100000110101001110100;
   assign mem[13081] = 32'b00000011001100010000010100010100;
   assign mem[13082] = 32'b00000011110000010001011111101100;
   assign mem[13083] = 32'b11111110010001100000010001010000;
   assign mem[13084] = 32'b11111110011000111010011111100000;
   assign mem[13085] = 32'b11111110111010101000100011100000;
   assign mem[13086] = 32'b00000001010100111001000101011000;
   assign mem[13087] = 32'b11111110011110110101010000001110;
   assign mem[13088] = 32'b11111001011010010001001011001000;
   assign mem[13089] = 32'b11111101111000001001010000101000;
   assign mem[13090] = 32'b11111000010100110100110001010000;
   assign mem[13091] = 32'b00000101101100010000110110010000;
   assign mem[13092] = 32'b11110100101010101100101010010000;
   assign mem[13093] = 32'b00001101000010001011101010000000;
   assign mem[13094] = 32'b11111001110001000101010101001000;
   assign mem[13095] = 32'b00000010001101100101000000111000;
   assign mem[13096] = 32'b11101010111110101001111111100000;
   assign mem[13097] = 32'b11111011010110000010111101110000;
   assign mem[13098] = 32'b11110001000000011100011111010000;
   assign mem[13099] = 32'b00000101010010100011101000100000;
   assign mem[13100] = 32'b00001001010100010000011100000000;
   assign mem[13101] = 32'b11111010011110001111011101010000;
   assign mem[13102] = 32'b11111111110000001010010101100010;
   assign mem[13103] = 32'b11111000011101110000100110010000;
   assign mem[13104] = 32'b11111010111111011010001001110000;
   assign mem[13105] = 32'b11111001100100111101000010100000;
   assign mem[13106] = 32'b11110111111010000001111001000000;
   assign mem[13107] = 32'b00000000101001000011010111001001;
   assign mem[13108] = 32'b11111111100011000011101101010101;
   assign mem[13109] = 32'b00000010001000011001011010001000;
   assign mem[13110] = 32'b11111111110010100011101011100101;
   assign mem[13111] = 32'b00000100110011011000111011111000;
   assign mem[13112] = 32'b11111111101010100000101001011100;
   assign mem[13113] = 32'b11111111010001101101010110010010;
   assign mem[13114] = 32'b11111110111001100011001011110000;
   assign mem[13115] = 32'b11111110011101101010100110101110;
   assign mem[13116] = 32'b11111010111101000011010111010000;
   assign mem[13117] = 32'b11110111000110110110101000010000;
   assign mem[13118] = 32'b00000011100111000010100111110000;
   assign mem[13119] = 32'b00000000001100000100101100010000;
   assign mem[13120] = 32'b00000100011010011101011011001000;
   assign mem[13121] = 32'b00001010110011100011110011110000;
   assign mem[13122] = 32'b00000001110010100110011100111100;
   assign mem[13123] = 32'b11110111010111011011010111010000;
   assign mem[13124] = 32'b00000100000011001101110010101000;
   assign mem[13125] = 32'b00000011001010111110101100110000;
   assign mem[13126] = 32'b11110100001100101011111001010000;
   assign mem[13127] = 32'b00000100010011111100011101111000;
   assign mem[13128] = 32'b00000100111110001101010010001000;
   assign mem[13129] = 32'b11110100111000100001011111100000;
   assign mem[13130] = 32'b00001100000101001000000010010000;
   assign mem[13131] = 32'b00000010100110001101110100101000;
   assign mem[13132] = 32'b00000001100110100000001010100110;
   assign mem[13133] = 32'b11110110111010111100000010100000;
   assign mem[13134] = 32'b11110110110110110011101000000000;
   assign mem[13135] = 32'b11110100101111110110011001010000;
   assign mem[13136] = 32'b11111110000001101001101100001100;
   assign mem[13137] = 32'b00001010001110110111111000010000;
   assign mem[13138] = 32'b11111110001001001101010000000100;
   assign mem[13139] = 32'b11111101011001110110110110100100;
   assign mem[13140] = 32'b00000011011011010001010110011100;
   assign mem[13141] = 32'b00000111000100110001011101001000;
   assign mem[13142] = 32'b00000000001100111011110011010111;
   assign mem[13143] = 32'b11111111101001110101101000010100;
   assign mem[13144] = 32'b11111110111110001010001001101110;
   assign mem[13145] = 32'b00000011011001110001000010001000;
   assign mem[13146] = 32'b00000001011010001100111111011100;
   assign mem[13147] = 32'b11111010000110101111110101110000;
   assign mem[13148] = 32'b00000010000011111000000110001100;
   assign mem[13149] = 32'b00000000100110100000101100100101;
   assign mem[13150] = 32'b11110000010110100100101100000000;
   assign mem[13151] = 32'b00000101101000011001000011001000;
   assign mem[13152] = 32'b00000100110110110100100111100000;
   assign mem[13153] = 32'b11111001010100110011110000110000;
   assign mem[13154] = 32'b00000010110010010011000010000100;
   assign mem[13155] = 32'b00000101101011000100111000000000;
   assign mem[13156] = 32'b11101111001010100100100001000000;
   assign mem[13157] = 32'b11111111010011110111111101101101;
   assign mem[13158] = 32'b11111010011100010000110001000000;
   assign mem[13159] = 32'b00000001000110001000100100100010;
   assign mem[13160] = 32'b00000001101000110011010110101110;
   assign mem[13161] = 32'b00000011001111000100111110010000;
   assign mem[13162] = 32'b11111110110110011110111111111110;
   assign mem[13163] = 32'b00000100010110000110001011101000;
   assign mem[13164] = 32'b11111111101000001101001101100101;
   assign mem[13165] = 32'b00000011011111000010101001000000;
   assign mem[13166] = 32'b11111011011011000101101001100000;
   assign mem[13167] = 32'b00000000010001001011101000001010;
   assign mem[13168] = 32'b11110000100000101010011000100000;
   assign mem[13169] = 32'b11111110001011001000111110000000;
   assign mem[13170] = 32'b11110101011010110011010111100000;
   assign mem[13171] = 32'b00000111101110010101101010111000;
   assign mem[13172] = 32'b11111110001100011111110100111010;
   assign mem[13173] = 32'b00000011100110111001001110011000;
   assign mem[13174] = 32'b00000000100001110011010110110100;
   assign mem[13175] = 32'b00000011110101110101000100111100;
   assign mem[13176] = 32'b11110101011010101110101000010000;
   assign mem[13177] = 32'b11111001000101101001001001101000;
   assign mem[13178] = 32'b11111010000000110111000001100000;
   assign mem[13179] = 32'b00000111100010010100010001011000;
   assign mem[13180] = 32'b11111110110101110110100111100100;
   assign mem[13181] = 32'b11111101101000011100001011110100;
   assign mem[13182] = 32'b00000010010100101100110001101000;
   assign mem[13183] = 32'b00000111001011011001101011101000;
   assign mem[13184] = 32'b00000110110001111101001011010000;
   assign mem[13185] = 32'b00000000001110000101100001101011;
   assign mem[13186] = 32'b11111011110101011101011010101000;
   assign mem[13187] = 32'b11110110101100101011010001000000;
   assign mem[13188] = 32'b11110111100101110000010101110000;
   assign mem[13189] = 32'b11111101111011100110100011011100;
   assign mem[13190] = 32'b11111101010010111111011000101000;
   assign mem[13191] = 32'b00001000100100011000010010000000;
   assign mem[13192] = 32'b11111100100000100010001000111100;
   assign mem[13193] = 32'b00000111111001111010101101101000;
   assign mem[13194] = 32'b00000100001001010101111101010000;
   assign mem[13195] = 32'b11111111111100001001111110110101;
   assign mem[13196] = 32'b11110101100110001101011010010000;
   assign mem[13197] = 32'b00000011001001111101110001110000;
   assign mem[13198] = 32'b11110100001000101010011010000000;
   assign mem[13199] = 32'b00000000010000100001001111100101;
   assign mem[13200] = 32'b00000000110110110100000010000111;
   assign mem[13201] = 32'b11101100011010110101010010100000;
   assign mem[13202] = 32'b00000001001100011000000001000000;
   assign mem[13203] = 32'b00000010010011111001100110110100;
   assign mem[13204] = 32'b00000000010001000000100101010110;
   assign mem[13205] = 32'b11111110110010101010000100100010;
   assign mem[13206] = 32'b00000000110001100011010111101111;
   assign mem[13207] = 32'b11110010100101111011011001000000;
   assign mem[13208] = 32'b00000100011111100010100001011000;
   assign mem[13209] = 32'b11111110111111110011000110100000;
   assign mem[13210] = 32'b00000010011010110110101101101000;
   assign mem[13211] = 32'b00000110100101011111000110110000;
   assign mem[13212] = 32'b11111110011101010000100101010000;
   assign mem[13213] = 32'b11111101011000111100101111010100;
   assign mem[13214] = 32'b00000001101110011111110010101110;
   assign mem[13215] = 32'b00000100011010000101011001010000;
   assign mem[13216] = 32'b00000010010000011000110101100000;
   assign mem[13217] = 32'b11111010110011010010011010100000;
   assign mem[13218] = 32'b11111000000111100101110111001000;
   assign mem[13219] = 32'b11111101110111100001101100110100;
   assign mem[13220] = 32'b00000001001101110010101110001100;
   assign mem[13221] = 32'b00000010100110001101010111000100;
   assign mem[13222] = 32'b00000000000100000010001100111100;
   assign mem[13223] = 32'b11111101010100111001001000011100;
   assign mem[13224] = 32'b00000010101011100110111011010000;
   assign mem[13225] = 32'b11111111011101111010000010111101;
   assign mem[13226] = 32'b11111111011100110100111010101001;
   assign mem[13227] = 32'b11111011001000010101100111101000;
   assign mem[13228] = 32'b00000010111010011110110000111100;
   assign mem[13229] = 32'b00000000011011001000010110101000;
   assign mem[13230] = 32'b11111110100011000111000000110000;
   assign mem[13231] = 32'b00000101100000011100101000010000;
   assign mem[13232] = 32'b00000110011110010100101001010000;
   assign mem[13233] = 32'b00000110100001110100010010010000;
   assign mem[13234] = 32'b00000011111101100010000010011000;
   assign mem[13235] = 32'b11110011111101000100100010010000;
   assign mem[13236] = 32'b00000011010001110010001100000000;
   assign mem[13237] = 32'b11111011100001111101100010101000;
   assign mem[13238] = 32'b11111101100111011011000011001000;
   assign mem[13239] = 32'b11111111011110011010100101111111;
   assign mem[13240] = 32'b00000001101011110101100110101000;
   assign mem[13241] = 32'b11110001100100001111010100000000;
   assign mem[13242] = 32'b11111110000011101011001110001100;
   assign mem[13243] = 32'b00000000000010100011100100001100;
   assign mem[13244] = 32'b11111110110100111101100101111010;
   assign mem[13245] = 32'b00000000100110001001010010001011;
   assign mem[13246] = 32'b00000000100010011011000111001010;
   assign mem[13247] = 32'b11111100100001100011000100010000;
   assign mem[13248] = 32'b00000100110000011010011010001000;
   assign mem[13249] = 32'b00000000010011010010000110001010;
   assign mem[13250] = 32'b11111101100101110000001101110100;
   assign mem[13251] = 32'b00000001101001110001011101100110;
   assign mem[13252] = 32'b00000000000101101111110001100111;
   assign mem[13253] = 32'b00000001111101100110100001000100;
   assign mem[13254] = 32'b11111010100111001111101100001000;
   assign mem[13255] = 32'b00000100010011000111001100110000;
   assign mem[13256] = 32'b11110111011000101000100101010000;
   assign mem[13257] = 32'b00000100011000011101011000101000;
   assign mem[13258] = 32'b00000000101011001101010010001110;
   assign mem[13259] = 32'b11111001101111010101111010011000;
   assign mem[13260] = 32'b00000110101100110110111101000000;
   assign mem[13261] = 32'b00000001110110010101101001111110;
   assign mem[13262] = 32'b00000111011111101000010100001000;
   assign mem[13263] = 32'b00000110011110100011000101101000;
   assign mem[13264] = 32'b11111110010000011111001110100100;
   assign mem[13265] = 32'b11111101000000010001110100011100;
   assign mem[13266] = 32'b00000010010100110010111100111000;
   assign mem[13267] = 32'b11110010111011011000010001000000;
   assign mem[13268] = 32'b00000001110000011111000111010110;
   assign mem[13269] = 32'b11111000011000001011111110000000;
   assign mem[13270] = 32'b11111111000101000101100001101010;
   assign mem[13271] = 32'b11111110011010010010111011111000;
   assign mem[13272] = 32'b00000001001111110111111011101100;
   assign mem[13273] = 32'b11111110100100110011111100010000;
   assign mem[13274] = 32'b11111101100110000111001001000000;
   assign mem[13275] = 32'b00000001100110100010100001001010;
   assign mem[13276] = 32'b00000000001001011011011111010001;
   assign mem[13277] = 32'b00000011011011001000011101100100;
   assign mem[13278] = 32'b11111110000011001110011001001100;
   assign mem[13279] = 32'b11111100100100010000111110001100;
   assign mem[13280] = 32'b00000010000011101011111110101000;
   assign mem[13281] = 32'b11111001010101111001010101110000;
   assign mem[13282] = 32'b00001000010011110100100100100000;
   assign mem[13283] = 32'b11111000010010111110000111111000;
   assign mem[13284] = 32'b00001000010011111100010001010000;
   assign mem[13285] = 32'b11111100100100000001100100011100;
   assign mem[13286] = 32'b00000000011001000100011110000011;
   assign mem[13287] = 32'b11111100000111011100101110111000;
   assign mem[13288] = 32'b11111001000111011101011010011000;
   assign mem[13289] = 32'b11111110000111111110101000000000;
   assign mem[13290] = 32'b11111001100111000011010010000000;
   assign mem[13291] = 32'b00000011011010011010101010110000;
   assign mem[13292] = 32'b00000011101011111011011111011100;
   assign mem[13293] = 32'b11111010110000011001110001011000;
   assign mem[13294] = 32'b11110011101111010011010010010000;
   assign mem[13295] = 32'b11110111100101100001001000110000;
   assign mem[13296] = 32'b11111100000000111010011100001000;
   assign mem[13297] = 32'b00001001111010100001001001100000;
   assign mem[13298] = 32'b00000000000011011110110000100110;
   assign mem[13299] = 32'b00000011100001111000111011111000;
   assign mem[13300] = 32'b00000011111111101101101001010100;
   assign mem[13301] = 32'b00000000111010101111101111001010;
   assign mem[13302] = 32'b11111110111111100100101000101000;
   assign mem[13303] = 32'b11110111101010001001001101110000;
   assign mem[13304] = 32'b11111011111011110111011001001000;
   assign mem[13305] = 32'b11111110011000101000001011101110;
   assign mem[13306] = 32'b11111110111100000111001111011010;
   assign mem[13307] = 32'b00000010111010101010001110110000;
   assign mem[13308] = 32'b11111011110001100001001110000000;
   assign mem[13309] = 32'b00000010011110110101110111000100;
   assign mem[13310] = 32'b00000010101100001010000100101100;
   assign mem[13311] = 32'b00000010010011100001110101010000;
   assign mem[13312] = 32'b00000000100001100001110110110111;
   assign mem[13313] = 32'b11111111010100111100001101100100;
   assign mem[13314] = 32'b11111101010101101110000010000000;
   assign mem[13315] = 32'b11111111101010101110111111101010;
   assign mem[13316] = 32'b11111111110100100100010110001001;
   assign mem[13317] = 32'b11110111010101100000011101000000;
   assign mem[13318] = 32'b00000001001111001100010001011100;
   assign mem[13319] = 32'b11111111001011100011110101011010;
   assign mem[13320] = 32'b00000001101011000001010101110010;
   assign mem[13321] = 32'b00000000000011011000000101010111;
   assign mem[13322] = 32'b00000100000111010100001000101000;
   assign mem[13323] = 32'b00000000000001010110100100100101;
   assign mem[13324] = 32'b00000000000010000100001100000111;
   assign mem[13325] = 32'b11111011011010001110111110011000;
   assign mem[13326] = 32'b11111010101011010010110000110000;
   assign mem[13327] = 32'b11110110010001110011100111100000;
   assign mem[13328] = 32'b00000010010011100110110001011100;
   assign mem[13329] = 32'b11111100001111100110010110100100;
   assign mem[13330] = 32'b11111101110110010001001011011000;
   assign mem[13331] = 32'b00001010010000010010001011010000;
   assign mem[13332] = 32'b11111011010111011000110111011000;
   assign mem[13333] = 32'b11111111101011010001110000100100;
   assign mem[13334] = 32'b00000011001001010100010011111000;
   assign mem[13335] = 32'b11111110101101101010111110010000;
   assign mem[13336] = 32'b11111111001000110001000000000011;
   assign mem[13337] = 32'b11111100101100000010011000101100;
   assign mem[13338] = 32'b00000010101000110101010000100000;
   assign mem[13339] = 32'b00000001000110110110010101011100;
   assign mem[13340] = 32'b00000010111111110010111111100000;
   assign mem[13341] = 32'b00000010001101001011001101100000;
   assign mem[13342] = 32'b00000010001000101001001101000000;
   assign mem[13343] = 32'b00000000011001001011111010100011;
   assign mem[13344] = 32'b11111110110011110001011000011010;
   assign mem[13345] = 32'b11111100110001100010010111100000;
   assign mem[13346] = 32'b11111110101101011000101101101000;
   assign mem[13347] = 32'b11110111010101011001011001110000;
   assign mem[13348] = 32'b00000110011001110110101101011000;
   assign mem[13349] = 32'b11111001010101110101100101111000;
   assign mem[13350] = 32'b11110110011100001001101101110000;
   assign mem[13351] = 32'b00010001111001011111111000100000;
   assign mem[13352] = 32'b00001001100111001001011111110000;
   assign mem[13353] = 32'b11111101111100111111010100010100;
   assign mem[13354] = 32'b00000011100001001111010000100100;
   assign mem[13355] = 32'b11111010110010100010110011000000;
   assign mem[13356] = 32'b11110000010101001000111111100000;
   assign mem[13357] = 32'b11111101000101000110100111100000;
   assign mem[13358] = 32'b00000001001010010000000011110110;
   assign mem[13359] = 32'b11110111011001010001111011100000;
   assign mem[13360] = 32'b00000010000101011100011100001100;
   assign mem[13361] = 32'b00000001100100101110101100001110;
   assign mem[13362] = 32'b00000011010011111111001111011100;
   assign mem[13363] = 32'b00000100011111000001001000010000;
   assign mem[13364] = 32'b11111010010010001011010010111000;
   assign mem[13365] = 32'b00000000100101101100000100100011;
   assign mem[13366] = 32'b11111110111011110000001101111000;
   assign mem[13367] = 32'b00000000100100111110001001001001;
   assign mem[13368] = 32'b11111011010111000100101000111000;
   assign mem[13369] = 32'b00000000111111001001011111010100;
   assign mem[13370] = 32'b00000001100101010101110110000000;
   assign mem[13371] = 32'b11111101000100011011000111100100;
   assign mem[13372] = 32'b00000001001110011101101101001010;
   assign mem[13373] = 32'b00000010011110001100010101001000;
   assign mem[13374] = 32'b11111011011011010011001001101000;
   assign mem[13375] = 32'b11111111101000011101110001111000;
   assign mem[13376] = 32'b11111110110100001100011100001000;
   assign mem[13377] = 32'b11110010001010100000111111010000;
   assign mem[13378] = 32'b11111111001010011110001011110001;
   assign mem[13379] = 32'b11111111110110011011111101011111;
   assign mem[13380] = 32'b11110000101001001111110000000000;
   assign mem[13381] = 32'b00000100000101011100100110101000;
   assign mem[13382] = 32'b11110001000110010101011010010000;
   assign mem[13383] = 32'b00001010100101110111111101000000;
   assign mem[13384] = 32'b11110111010000101101100101010000;
   assign mem[13385] = 32'b00001000111001101000011001000000;
   assign mem[13386] = 32'b11110011000111101111001010010000;
   assign mem[13387] = 32'b00000010010000011111101110001000;
   assign mem[13388] = 32'b11110000000110011000111110010000;
   assign mem[13389] = 32'b00000101111010100010001000001000;
   assign mem[13390] = 32'b11111001000001001111000100110000;
   assign mem[13391] = 32'b11111111100010110011001001001100;
   assign mem[13392] = 32'b11111100000101100110100011010000;
   assign mem[13393] = 32'b00000100111011001111111110000000;
   assign mem[13394] = 32'b11111110011101011100100110001110;
   assign mem[13395] = 32'b00000001101010110001111011111010;
   assign mem[13396] = 32'b11110001101100011101101100000000;
   assign mem[13397] = 32'b00000001011011010111011100011100;
   assign mem[13398] = 32'b00000000111101110111010001011000;
   assign mem[13399] = 32'b00000110111101010110011111010000;
   assign mem[13400] = 32'b11100001000101111100001001000000;
   assign mem[13401] = 32'b00000101101000001101111100110000;
   assign mem[13402] = 32'b11111010110010100010001110010000;
   assign mem[13403] = 32'b00000011110110101111000011111100;
   assign mem[13404] = 32'b11111111011001100101111101101011;
   assign mem[13405] = 32'b00000101100100101000111011101000;
   assign mem[13406] = 32'b11101000010100101000010111000000;
   assign mem[13407] = 32'b00000001001110101101000101111110;
   assign mem[13408] = 32'b11111011010001000010011010110000;
   assign mem[13409] = 32'b00000101010101101111111111100000;
   assign mem[13410] = 32'b00000011011110111011111001001000;
   assign mem[13411] = 32'b00000000010100011000111111110011;
   assign mem[13412] = 32'b00000010001000010100110001011000;
   assign mem[13413] = 32'b11101111011110110111101101000000;
   assign mem[13414] = 32'b11111111010111000010101110010100;
   assign mem[13415] = 32'b11110100110000101010010010110000;
   assign mem[13416] = 32'b11110111111100001000010000000000;
   assign mem[13417] = 32'b00001000001010101111011000000000;
   assign mem[13418] = 32'b00000011011001000110001110110000;
   assign mem[13419] = 32'b11111111000101111101011010011101;
   assign mem[13420] = 32'b00000111010100100100100010110000;
   assign mem[13421] = 32'b00000010100011010100000011000100;
   assign mem[13422] = 32'b00000110100001011010010011001000;
   assign mem[13423] = 32'b00000010101100111000110000001000;
   assign mem[13424] = 32'b11111000100010001011011111011000;
   assign mem[13425] = 32'b11111011010000010011101111111000;
   assign mem[13426] = 32'b11111111011111000000000101011110;
   assign mem[13427] = 32'b00000000010101110011111001100010;
   assign mem[13428] = 32'b11111111100011100100101000000011;
   assign mem[13429] = 32'b11111011000001100111100000110000;
   assign mem[13430] = 32'b00000010000111001010110101000000;
   assign mem[13431] = 32'b00001011010001011100001011000000;
   assign mem[13432] = 32'b00000101001000100011000001000000;
   assign mem[13433] = 32'b11111101010101101011001011100000;
   assign mem[13434] = 32'b11110111110000001110000000100000;
   assign mem[13435] = 32'b11111001000111101111011000100000;
   assign mem[13436] = 32'b11111110011110100011100100100110;
   assign mem[13437] = 32'b11111010110011011010100000000000;
   assign mem[13438] = 32'b00000000001101100100011000101000;
   assign mem[13439] = 32'b11111100101111101100000100010100;
   assign mem[13440] = 32'b00000001001011111100110100101010;
   assign mem[13441] = 32'b11111011100001111101111001011000;
   assign mem[13442] = 32'b11111110101001100011100101001010;
   assign mem[13443] = 32'b00000010010001101011010110111000;
   assign mem[13444] = 32'b11111101011111111011011010110000;
   assign mem[13445] = 32'b11111111001101110010101111111100;
   assign mem[13446] = 32'b11111110000111001100010010111100;
   assign mem[13447] = 32'b11110110001111010111000000110000;
   assign mem[13448] = 32'b00000011100001110001111010011100;
   assign mem[13449] = 32'b11111101001001100000010101100000;
   assign mem[13450] = 32'b00001011011011001110011100100000;
   assign mem[13451] = 32'b11111100001011001001100001001000;
   assign mem[13452] = 32'b11110101001001011111011101100000;
   assign mem[13453] = 32'b00000010111010001011000110000000;
   assign mem[13454] = 32'b11110100011110011101100111010000;
   assign mem[13455] = 32'b00000010011101001000010010000100;
   assign mem[13456] = 32'b11111110001001110101001010011000;
   assign mem[13457] = 32'b00000101000100001001011100010000;
   assign mem[13458] = 32'b11110101001011110100000100000000;
   assign mem[13459] = 32'b00000110000011111001001100001000;
   assign mem[13460] = 32'b11111110010010110010000000000010;
   assign mem[13461] = 32'b11110101101011101111011011000000;
   assign mem[13462] = 32'b00000011001100001100011011101100;
   assign mem[13463] = 32'b00000010111001011101001001111000;
   assign mem[13464] = 32'b11111111100010001010100110000101;
   assign mem[13465] = 32'b00000010101000100001011110110100;
   assign mem[13466] = 32'b00000100100110000111101101111000;
   assign mem[13467] = 32'b11100010110001111011001111000000;
   assign mem[13468] = 32'b00000110011000011110011101011000;
   assign mem[13469] = 32'b11111101001110010000100100111100;
   assign mem[13470] = 32'b00000000110110101010101010111001;
   assign mem[13471] = 32'b11111101100101010101011100110000;
   assign mem[13472] = 32'b11111100101001101001010100110000;
   assign mem[13473] = 32'b00000010001001100001011100101000;
   assign mem[13474] = 32'b11111100001111010101011000110100;
   assign mem[13475] = 32'b00000100010010010011001000010000;
   assign mem[13476] = 32'b00000001110000010010100000000110;
   assign mem[13477] = 32'b00000000101111100111101000111011;
   assign mem[13478] = 32'b11111011111100100000101011010000;
   assign mem[13479] = 32'b00000100110000001111000110110000;
   assign mem[13480] = 32'b11111111000101001001000100000110;
   assign mem[13481] = 32'b00000000110110000001001010111110;
   assign mem[13482] = 32'b00000010101011011001001111110000;
   assign mem[13483] = 32'b11111111011101110001001000100000;
   assign mem[13484] = 32'b11111110110000000111111101111110;
   assign mem[13485] = 32'b00000011111010010111000001000000;
   assign mem[13486] = 32'b11111100000011011100111011111100;
   assign mem[13487] = 32'b00000000011111011110111110110101;
   assign mem[13488] = 32'b11110111001100111001001111010000;
   assign mem[13489] = 32'b00000101010001111000100000001000;
   assign mem[13490] = 32'b00000000011011010000111010100110;
   assign mem[13491] = 32'b11111110111010100110011111100010;
   assign mem[13492] = 32'b11111111011001111100101011010111;
   assign mem[13493] = 32'b11110101110101010001011000010000;
   assign mem[13494] = 32'b00000100001000001100110011100000;
   assign mem[13495] = 32'b11110111111110011010001011110000;
   assign mem[13496] = 32'b11111010111110011000011010101000;
   assign mem[13497] = 32'b00000110111010101010000001011000;
   assign mem[13498] = 32'b00000011101011000111111111101000;
   assign mem[13499] = 32'b00000000010010111011010010010101;
   assign mem[13500] = 32'b11101111101110001011000011100000;
   assign mem[13501] = 32'b00001111000011111100000000110000;
   assign mem[13502] = 32'b00001010110011001110010101100000;
   assign mem[13503] = 32'b11110011110111010110100011110000;
   assign mem[13504] = 32'b11111110000100001010100011001100;
   assign mem[13505] = 32'b00000000011000000111111000001110;
   assign mem[13506] = 32'b11100110000110101100101111000000;
   assign mem[13507] = 32'b00001101100110000101011011010000;
   assign mem[13508] = 32'b11111101001001110001011010100000;
   assign mem[13509] = 32'b11111010000011010101000101101000;
   assign mem[13510] = 32'b11110110011011011111101111100000;
   assign mem[13511] = 32'b00000101110000110111110001101000;
   assign mem[13512] = 32'b11111100110111010101111110101000;
   assign mem[13513] = 32'b11110111100010000100111000000000;
   assign mem[13514] = 32'b00000010001001111100001010100000;
   assign mem[13515] = 32'b11111100110101011110111110110000;
   assign mem[13516] = 32'b11111001111100110101000101000000;
   assign mem[13517] = 32'b00000101011111000110000001110000;
   assign mem[13518] = 32'b11110110000100111111010000010000;
   assign mem[13519] = 32'b00000011101101011101110110100100;
   assign mem[13520] = 32'b11111110000101000111101111111100;
   assign mem[13521] = 32'b00000110111111000111001111011000;
   assign mem[13522] = 32'b11101100101010100110010111000000;
   assign mem[13523] = 32'b00001001000011011100010111000000;
   assign mem[13524] = 32'b11110101000101101100001001000000;
   assign mem[13525] = 32'b00001001111001110110101111100000;
   assign mem[13526] = 32'b11110010100000001101011100110000;
   assign mem[13527] = 32'b11110101110001111100001100100000;
   assign mem[13528] = 32'b11110000001110111011011000110000;
   assign mem[13529] = 32'b00000011011111000100111001001000;
   assign mem[13530] = 32'b11111111010110101110011011000001;
   assign mem[13531] = 32'b00000101001010100111001100111000;
   assign mem[13532] = 32'b00000101101010010000000110100000;
   assign mem[13533] = 32'b11110000100010001010000000100000;
   assign mem[13534] = 32'b00000000000001010100100111101000;
   assign mem[13535] = 32'b11101100111101010010100100000000;
   assign mem[13536] = 32'b11111001010101001001011101110000;
   assign mem[13537] = 32'b00000001011100110110001001110110;
   assign mem[13538] = 32'b00000011000011011010110110011000;
   assign mem[13539] = 32'b11111110100010111010101110010100;
   assign mem[13540] = 32'b00000010000101111101100100100000;
   assign mem[13541] = 32'b00001001001101110100111100010000;
   assign mem[13542] = 32'b11111001100001100001101010111000;
   assign mem[13543] = 32'b11111111111011010000100010000011;
   assign mem[13544] = 32'b00000010001100110110100111001000;
   assign mem[13545] = 32'b00001000100100110011110110000000;
   assign mem[13546] = 32'b11111001000010011110011010111000;
   assign mem[13547] = 32'b11111001100001000000000110000000;
   assign mem[13548] = 32'b11111100011000100101100010110100;
   assign mem[13549] = 32'b00000011111000001000110111010000;
   assign mem[13550] = 32'b11111110110101010011001011010010;
   assign mem[13551] = 32'b11111100011100011011101001010100;
   assign mem[13552] = 32'b11111101010001001001111001001000;
   assign mem[13553] = 32'b11111110100101101010010111011110;
   assign mem[13554] = 32'b11111001101011001011100011010000;
   assign mem[13555] = 32'b00000001101001110111100101111100;
   assign mem[13556] = 32'b00000011100111010011101000010100;
   assign mem[13557] = 32'b11111000000101100110010110011000;
   assign mem[13558] = 32'b00000000010110010101010001110101;
   assign mem[13559] = 32'b11111110101101011111101011010010;
   assign mem[13560] = 32'b00000111000000100101000000110000;
   assign mem[13561] = 32'b00000011011110001111000010011000;
   assign mem[13562] = 32'b11111110011000000101011011000110;
   assign mem[13563] = 32'b00000000110011101010110110100111;
   assign mem[13564] = 32'b11111000000110001110001111001000;
   assign mem[13565] = 32'b11111111110101001010010111110100;
   assign mem[13566] = 32'b00000010110101010101011010101100;
   assign mem[13567] = 32'b11100111010100001101011001100000;
   assign mem[13568] = 32'b00000110111000100011010111100000;
   assign mem[13569] = 32'b11111100010011100111101011010100;
   assign mem[13570] = 32'b11111010110001100010010110001000;
   assign mem[13571] = 32'b00001100111101111010101000000000;
   assign mem[13572] = 32'b11110111101011111010010001110000;
   assign mem[13573] = 32'b00000100000011100110110100000000;
   assign mem[13574] = 32'b11110001111101001000011011100000;
   assign mem[13575] = 32'b00000010111101001101110000001000;
   assign mem[13576] = 32'b11110110011110110010011100000000;
   assign mem[13577] = 32'b11100011111001000001000111000000;
   assign mem[13578] = 32'b00000100100011000110110111000000;
   assign mem[13579] = 32'b00000011100000000100011001011000;
   assign mem[13580] = 32'b00000001100111100101110010100010;
   assign mem[13581] = 32'b11111000011000010010011000111000;
   assign mem[13582] = 32'b00000010111101000101110111101100;
   assign mem[13583] = 32'b11111111010101111110111100110000;
   assign mem[13584] = 32'b11110101111100001111000101000000;
   assign mem[13585] = 32'b00000000101100111010110101101011;
   assign mem[13586] = 32'b11111101101110100110100110111100;
   assign mem[13587] = 32'b11110100101100001101101010000000;
   assign mem[13588] = 32'b00000101010111001101101100100000;
   assign mem[13589] = 32'b11111010010100001011001100111000;
   assign mem[13590] = 32'b11111001010011010100110000101000;
   assign mem[13591] = 32'b00000100100011101011110010010000;
   assign mem[13592] = 32'b11111010011110100110000111111000;
   assign mem[13593] = 32'b11111000011110111001100101000000;
   assign mem[13594] = 32'b00000001101011101000001101100100;
   assign mem[13595] = 32'b11111101111111000100100100101100;
   assign mem[13596] = 32'b11111010101010010100010001001000;
   assign mem[13597] = 32'b00000001110001101111101100101100;
   assign mem[13598] = 32'b00000010111111110000010100101100;
   assign mem[13599] = 32'b00000010010111010011100010010000;
   assign mem[13600] = 32'b00000101110100101110110100001000;
   assign mem[13601] = 32'b11111100101011000000001100010000;
   assign mem[13602] = 32'b00000011110001010110011000101000;
   assign mem[13603] = 32'b00000001011010111101110010110000;
   assign mem[13604] = 32'b11111011001110001111101100001000;
   assign mem[13605] = 32'b00000001101110000001110000000100;
   assign mem[13606] = 32'b00000010110101101100011000011100;
   assign mem[13607] = 32'b11110110000000100011110010010000;
   assign mem[13608] = 32'b00000001111101111100100010100110;
   assign mem[13609] = 32'b11111011101111110110111010011000;
   assign mem[13610] = 32'b00000100100111000111010011000000;
   assign mem[13611] = 32'b11111111000000101100000101100100;
   assign mem[13612] = 32'b11111111011111101110111011111001;
   assign mem[13613] = 32'b11111101101110010000101010100100;
   assign mem[13614] = 32'b11110100010010110101101010100000;
   assign mem[13615] = 32'b00000001100010001010001111111110;
   assign mem[13616] = 32'b00000001101101011111011001010110;
   assign mem[13617] = 32'b00000000101010010001100000011110;
   assign mem[13618] = 32'b00000010111110010100000110110100;
   assign mem[13619] = 32'b11110100010100010111110100010000;
   assign mem[13620] = 32'b00000100110110100001111001110000;
   assign mem[13621] = 32'b00000010110000001000110100110100;
   assign mem[13622] = 32'b00000101010010001010111001110000;
   assign mem[13623] = 32'b11111101001100101111101000011000;
   assign mem[13624] = 32'b00000000100100000101010010010110;
   assign mem[13625] = 32'b11111101110000001011100000010100;
   assign mem[13626] = 32'b11111100001001111110010001101100;
   assign mem[13627] = 32'b11111010111101010101001011011000;
   assign mem[13628] = 32'b11111110000110110110011001000100;
   assign mem[13629] = 32'b11111100001101101101110110110100;
   assign mem[13630] = 32'b00000111100110010010001001101000;
   assign mem[13631] = 32'b00000101011011001011011010111000;
   assign mem[13632] = 32'b11111100001010001011001111100000;
   assign mem[13633] = 32'b00000100110011010100000100011000;
   assign mem[13634] = 32'b00000010001000010110011011111100;
   assign mem[13635] = 32'b00000100100100111010000000011000;
   assign mem[13636] = 32'b11100111010100111111010010000000;
   assign mem[13637] = 32'b11111111000001000001110001010111;
   assign mem[13638] = 32'b00000000001011101010100010101111;
   assign mem[13639] = 32'b11111100001001001000100001001000;
   assign mem[13640] = 32'b00000101001010100001100001011000;
   assign mem[13641] = 32'b00000010101000110010110000100000;
   assign mem[13642] = 32'b00000001001001000110000010110100;
   assign mem[13643] = 32'b11101101111101010000110001000000;
   assign mem[13644] = 32'b11111111000110010011100100110100;
   assign mem[13645] = 32'b11110110010100011001101100100000;
   assign mem[13646] = 32'b00000000110010011101111000011001;
   assign mem[13647] = 32'b00000010101000010011000111111100;
   assign mem[13648] = 32'b00000010100110110010000101111000;
   assign mem[13649] = 32'b11110110001111011110101100110000;
   assign mem[13650] = 32'b11111101011111101001101000011000;
   assign mem[13651] = 32'b00000001111111010100011011101110;
   assign mem[13652] = 32'b11111011001001100110000011011000;
   assign mem[13653] = 32'b00001000001001111011011011100000;
   assign mem[13654] = 32'b11111010100110101110000100011000;
   assign mem[13655] = 32'b00000101100101010110100111010000;
   assign mem[13656] = 32'b11110110010011011011100100010000;
   assign mem[13657] = 32'b11111000100010001111101110101000;
   assign mem[13658] = 32'b11111011011011101111001101001000;
   assign mem[13659] = 32'b00000000001010010010101011100000;
   assign mem[13660] = 32'b11111010100101110100111100100000;
   assign mem[13661] = 32'b00000100101000101001011100111000;
   assign mem[13662] = 32'b11111000011100000101010111100000;
   assign mem[13663] = 32'b11110110100001110011001101010000;
   assign mem[13664] = 32'b00001001001001000111101011110000;
   assign mem[13665] = 32'b00000111000010011111111101101000;
   assign mem[13666] = 32'b11110110010000111101011010100000;
   assign mem[13667] = 32'b00000110001001111010100000101000;
   assign mem[13668] = 32'b11111000110100101001011101001000;
   assign mem[13669] = 32'b00000111001110100011110111110000;
   assign mem[13670] = 32'b00000010000111001110001001111000;
   assign mem[13671] = 32'b11111010000101110010000001001000;
   assign mem[13672] = 32'b00000001111010111110000011011110;
   assign mem[13673] = 32'b11111111110000111110001111101100;
   assign mem[13674] = 32'b11110110010011011010011100010000;
   assign mem[13675] = 32'b11111110110001010100110111011010;
   assign mem[13676] = 32'b00000010001010010111101011011100;
   assign mem[13677] = 32'b11110011100001000110000100110000;
   assign mem[13678] = 32'b00000011000011110100100101100000;
   assign mem[13679] = 32'b11110110000111111010101011010000;
   assign mem[13680] = 32'b00000010011000011111100011001100;
   assign mem[13681] = 32'b11110001001110100100011100010000;
   assign mem[13682] = 32'b00000100100000110011101100011000;
   assign mem[13683] = 32'b11111111111111000001000011011010;
   assign mem[13684] = 32'b11110101001110110001001001000000;
   assign mem[13685] = 32'b00000011110111000101000101111000;
   assign mem[13686] = 32'b00000010000101100000001010101100;
   assign mem[13687] = 32'b11110000001010100010001100000000;
   assign mem[13688] = 32'b00000110011001010110111101010000;
   assign mem[13689] = 32'b11111000110011101101111111001000;
   assign mem[13690] = 32'b11111101111010001011001101000000;
   assign mem[13691] = 32'b00010111000101101101001001100000;
   assign mem[13692] = 32'b00000011010011111010010000101000;
   assign mem[13693] = 32'b11111000011011111100111011010000;
   assign mem[13694] = 32'b00000001011100001001100100001110;
   assign mem[13695] = 32'b00001001101111101001001011110000;
   assign mem[13696] = 32'b11110011000000000110111001000000;
   assign mem[13697] = 32'b00001010110010100110100000110000;
   assign mem[13698] = 32'b11111110001001010100010100011000;
   assign mem[13699] = 32'b11110010110101100100101000100000;
   assign mem[13700] = 32'b00001011000001110011101101010000;
   assign mem[13701] = 32'b11111101100010101100101111101000;
   assign mem[13702] = 32'b00000000110100100001001011101111;
   assign mem[13703] = 32'b11111010011001110101011101011000;
   assign mem[13704] = 32'b11111011110100100010010001010000;
   assign mem[13705] = 32'b11111111110101110010011001100110;
   assign mem[13706] = 32'b00000100010011110111110000011000;
   assign mem[13707] = 32'b11111011101010100110111000010000;
   assign mem[13708] = 32'b00001000111110011000001110000000;
   assign mem[13709] = 32'b11101011110100011010010101000000;
   assign mem[13710] = 32'b11100110011111000000011011100000;
   assign mem[13711] = 32'b00000100010100111001110111100000;
   assign mem[13712] = 32'b00000011001111000110111111110100;
   assign mem[13713] = 32'b00000110111111111001000100001000;
   assign mem[13714] = 32'b11111110010111001000101101110110;
   assign mem[13715] = 32'b00001001111101111111001011010000;
   assign mem[13716] = 32'b11101100100110111111100111100000;
   assign mem[13717] = 32'b00000000001101100111010101011000;
   assign mem[13718] = 32'b11111001100011011000110110100000;
   assign mem[13719] = 32'b00000100000111111011101010010000;
   assign mem[13720] = 32'b00000001101000111001010001111100;
   assign mem[13721] = 32'b00000101000111010011011000100000;
   assign mem[13722] = 32'b00000000010011111110110010100011;
   assign mem[13723] = 32'b11111101011110011111100001000000;
   assign mem[13724] = 32'b11111010110010101101110111100000;
   assign mem[13725] = 32'b11111100110100100101101100010100;
   assign mem[13726] = 32'b00000001011111101010110000000110;
   assign mem[13727] = 32'b11110111010110100011101011000000;
   assign mem[13728] = 32'b00000010010101101000010001110100;
   assign mem[13729] = 32'b00000001111111101101111000000100;
   assign mem[13730] = 32'b11111010101110000100110100100000;
   assign mem[13731] = 32'b00001101100101100000110001010000;
   assign mem[13732] = 32'b11110011110000100010011011110000;
   assign mem[13733] = 32'b00001000100001111101000011100000;
   assign mem[13734] = 32'b11110000111010000111111001010000;
   assign mem[13735] = 32'b00001011100100011010010000010000;
   assign mem[13736] = 32'b11101111010000011100100000000000;
   assign mem[13737] = 32'b11110111100100000001010100000000;
   assign mem[13738] = 32'b11101111010011001011101001100000;
   assign mem[13739] = 32'b00000110101100101010001110111000;
   assign mem[13740] = 32'b00000011111101100101001001001000;
   assign mem[13741] = 32'b00010110000000001101010101000000;
   assign mem[13742] = 32'b11111001000100111110100000000000;
   assign mem[13743] = 32'b11110011101110110011011011100000;
   assign mem[13744] = 32'b00000100101111000111000100101000;
   assign mem[13745] = 32'b11111001110000101000100001010000;
   assign mem[13746] = 32'b00000000011010000111001110101111;
   assign mem[13747] = 32'b00000011100001101101110101011100;
   assign mem[13748] = 32'b00000001010111010001111111111110;
   assign mem[13749] = 32'b11111011100011111110000100011000;
   assign mem[13750] = 32'b11111110100100001111100111101110;
   assign mem[13751] = 32'b11111111010010011101101011011011;
   assign mem[13752] = 32'b00000000001100110101001101101101;
   assign mem[13753] = 32'b00000001100100001101010010111000;
   assign mem[13754] = 32'b11111110010010111010100101010000;
   assign mem[13755] = 32'b00000010001010101011110001111100;
   assign mem[13756] = 32'b00000000111000101000100111110000;
   assign mem[13757] = 32'b11111000100101111010110111010000;
   assign mem[13758] = 32'b11111111011011001111001110101100;
   assign mem[13759] = 32'b00000000101001010100110101100101;
   assign mem[13760] = 32'b11111100001011101111111011000000;
   assign mem[13761] = 32'b11111111011011001111000000110011;
   assign mem[13762] = 32'b00000010101101000001110010111100;
   assign mem[13763] = 32'b11111011101011010011100001010000;
   assign mem[13764] = 32'b00000111001101101001011101011000;
   assign mem[13765] = 32'b00000010010011000100100011100000;
   assign mem[13766] = 32'b11110110101010010100001011100000;
   assign mem[13767] = 32'b00000101001110011100100010111000;
   assign mem[13768] = 32'b00000100110101010001110101111000;
   assign mem[13769] = 32'b00000110010001010010001010010000;
   assign mem[13770] = 32'b11111000101110010011001011110000;
   assign mem[13771] = 32'b00000111000111011000101110101000;
   assign mem[13772] = 32'b11111011110000011000111110010000;
   assign mem[13773] = 32'b11110101010100000110100011110000;
   assign mem[13774] = 32'b00001000111011001010110100100000;
   assign mem[13775] = 32'b11110011100100111000101101100000;
   assign mem[13776] = 32'b11111010110000000001011110010000;
   assign mem[13777] = 32'b00000101101000110000010101011000;
   assign mem[13778] = 32'b11111100101100101001110101101000;
   assign mem[13779] = 32'b00000100011100001111110011010000;
   assign mem[13780] = 32'b00000010011100011101000011100000;
   assign mem[13781] = 32'b00000001011101100110100011110010;
   assign mem[13782] = 32'b11111110010001101010100010101110;
   assign mem[13783] = 32'b11111110001001100101001111100000;
   assign mem[13784] = 32'b11111111101000011101101101111000;
   assign mem[13785] = 32'b00000000011111010011011100000000;
   assign mem[13786] = 32'b00000000010111100110001000001100;
   assign mem[13787] = 32'b11111001111011111010001111110000;
   assign mem[13788] = 32'b11111110000100000011000101101110;
   assign mem[13789] = 32'b11111111101001101010110110001000;
   assign mem[13790] = 32'b11101100011011010110111100000000;
   assign mem[13791] = 32'b00001101110110100010011101000000;
   assign mem[13792] = 32'b00000110011011010101110110001000;
   assign mem[13793] = 32'b00001010011010110110100010100000;
   assign mem[13794] = 32'b11111011011100111101101010101000;
   assign mem[13795] = 32'b00000111010011010011000100011000;
   assign mem[13796] = 32'b11101110000111100000011001100000;
   assign mem[13797] = 32'b00001001010111011001110110010000;
   assign mem[13798] = 32'b11101101110010011010101100100000;
   assign mem[13799] = 32'b11111010110110111110011000010000;
   assign mem[13800] = 32'b11111111000010001010011010001010;
   assign mem[13801] = 32'b11111010011100000010110010000000;
   assign mem[13802] = 32'b00000000101000011000011110101010;
   assign mem[13803] = 32'b11111100101001000101101100001100;
   assign mem[13804] = 32'b11111001100110111010111111001000;
   assign mem[13805] = 32'b00000010110100111011001100111100;
   assign mem[13806] = 32'b11111001100001001111001011110000;
   assign mem[13807] = 32'b11111001011001000111100110001000;
   assign mem[13808] = 32'b11111101101100110101001100100100;
   assign mem[13809] = 32'b11111111101010100100010111100111;
   assign mem[13810] = 32'b00000011100001101110100010111000;
   assign mem[13811] = 32'b00001001110010001110010011010000;
   assign mem[13812] = 32'b11111110111000100100011010110110;
   assign mem[13813] = 32'b00000011000110011000010000110000;
   assign mem[13814] = 32'b11111010011111110100010011111000;
   assign mem[13815] = 32'b00000101110111111000101101100000;
   assign mem[13816] = 32'b11110010101000110001011000000000;
   assign mem[13817] = 32'b11110000111000001100111001100000;
   assign mem[13818] = 32'b11111100010100110101101100111100;
   assign mem[13819] = 32'b00000010000101010111011011010000;
   assign mem[13820] = 32'b00000010001100010110111010011000;
   assign mem[13821] = 32'b11111100001001000001101000110100;
   assign mem[13822] = 32'b00000000010011100000110101000101;
   assign mem[13823] = 32'b11111111101101100011100100110100;
   assign mem[13824] = 32'b11110111101110111001111011110000;
   assign mem[13825] = 32'b11111111110000000111111100010100;
   assign mem[13826] = 32'b11111110110001011001010000001100;
   assign mem[13827] = 32'b11111000001111010110110010101000;
   assign mem[13828] = 32'b00000010110011100011010101000100;
   assign mem[13829] = 32'b00000100000100000100001111100000;
   assign mem[13830] = 32'b11110101100101110000110010010000;
   assign mem[13831] = 32'b11111100001000100101000001100100;
   assign mem[13832] = 32'b00000010001000111111110010100100;
   assign mem[13833] = 32'b00000100100110000101000101011000;
   assign mem[13834] = 32'b11111111010011110010001101101101;
   assign mem[13835] = 32'b00001010110011100100000111100000;
   assign mem[13836] = 32'b11110101011011100110010111000000;
   assign mem[13837] = 32'b11111111011000011101001001111010;
   assign mem[13838] = 32'b11110001110111000101101011100000;
   assign mem[13839] = 32'b00000011000010000100100100010100;
   assign mem[13840] = 32'b00000101010010110000101101011000;
   assign mem[13841] = 32'b11110110010111001101101011100000;
   assign mem[13842] = 32'b00000011000100110011111100110000;
   assign mem[13843] = 32'b11111110111001000101000000001110;
   assign mem[13844] = 32'b11111000100101001000100001110000;
   assign mem[13845] = 32'b11111111101011001010000110010100;
   assign mem[13846] = 32'b00000101101110110100100011001000;
   assign mem[13847] = 32'b11111101011110100110010101010100;
   assign mem[13848] = 32'b00000001100101100001001111110010;
   assign mem[13849] = 32'b11111111001000100100101110000011;
   assign mem[13850] = 32'b00000000001111011011011110100110;
   assign mem[13851] = 32'b11111101111100110100110011000000;
   assign mem[13852] = 32'b00000011001011111111101011000100;
   assign mem[13853] = 32'b11111111100100001101111001111111;
   assign mem[13854] = 32'b11111011110101100100000001011000;
   assign mem[13855] = 32'b00000001001011111001001001001100;
   assign mem[13856] = 32'b00000000101101100011000101000111;
   assign mem[13857] = 32'b11111011000110100110111010001000;
   assign mem[13858] = 32'b11111010001000111110000010100000;
   assign mem[13859] = 32'b00000001001101001011011111000100;
   assign mem[13860] = 32'b11111111010011100111011011010101;
   assign mem[13861] = 32'b11111011110111001100010110101000;
   assign mem[13862] = 32'b11111110010110101100111000010000;
   assign mem[13863] = 32'b11111110101101000101111011110010;
   assign mem[13864] = 32'b11111101011011011001001101001100;
   assign mem[13865] = 32'b00000010000101111001101001111100;
   assign mem[13866] = 32'b00000010110110000001011111000000;
   assign mem[13867] = 32'b11111101110011111011110010010000;
   assign mem[13868] = 32'b11111100111101001010011011100000;
   assign mem[13869] = 32'b00000010101011100000000110000100;
   assign mem[13870] = 32'b00001001111011001101111101110000;
   assign mem[13871] = 32'b11111010100110100000010011110000;
   assign mem[13872] = 32'b00000111101001100110111101010000;
   assign mem[13873] = 32'b00000000011010111010110000100011;
   assign mem[13874] = 32'b11110111110010011111000110110000;
   assign mem[13875] = 32'b00000011001011111011000001010100;
   assign mem[13876] = 32'b11111111001010001011011111011000;
   assign mem[13877] = 32'b11110101010011000001101111010000;
   assign mem[13878] = 32'b11111001000011100010111111100000;
   assign mem[13879] = 32'b11111011011000011110111010011000;
   assign mem[13880] = 32'b00000010111101111100000100110100;
   assign mem[13881] = 32'b11111011111101110011100000110000;
   assign mem[13882] = 32'b00000100000001101111001110101000;
   assign mem[13883] = 32'b11111111110001111100000100010111;
   assign mem[13884] = 32'b11111001110111011110111111100000;
   assign mem[13885] = 32'b11111101010010011101100011010000;
   assign mem[13886] = 32'b00000011000110010111101010011000;
   assign mem[13887] = 32'b11101110010010000010011110000000;
   assign mem[13888] = 32'b00000101010000000101111000011000;
   assign mem[13889] = 32'b11111100011111100110010100101100;
   assign mem[13890] = 32'b00001011001000110011101100000000;
   assign mem[13891] = 32'b11110011010111111110101001010000;
   assign mem[13892] = 32'b11111111011000101010101100101111;
   assign mem[13893] = 32'b00000011100010110101010111011100;
   assign mem[13894] = 32'b00000100001001100011001101010000;
   assign mem[13895] = 32'b00000101100001001011100000011000;
   assign mem[13896] = 32'b11111010110001000100001100011000;
   assign mem[13897] = 32'b00000011000101001110110110111100;
   assign mem[13898] = 32'b11111101011000001001110001001000;
   assign mem[13899] = 32'b11111001100110000110001001111000;
   assign mem[13900] = 32'b00000101010001011000011100010000;
   assign mem[13901] = 32'b00000101011111100001010000000000;
   assign mem[13902] = 32'b11111011001011110101011101010000;
   assign mem[13903] = 32'b11110101010001110000110110100000;
   assign mem[13904] = 32'b11111110101010000101110111101000;
   assign mem[13905] = 32'b11111011010111100110000000110000;
   assign mem[13906] = 32'b00000101111111000100011100111000;
   assign mem[13907] = 32'b00000100010111100011000101010000;
   assign mem[13908] = 32'b00000010011010111000101110101000;
   assign mem[13909] = 32'b11111011110100111101001011100000;
   assign mem[13910] = 32'b00000010111110011001001000000100;
   assign mem[13911] = 32'b11111110010001101011010011010000;
   assign mem[13912] = 32'b00000010111110110000010100100000;
   assign mem[13913] = 32'b11111110101111001100001100101110;
   assign mem[13914] = 32'b11111101000011100101101110101100;
   assign mem[13915] = 32'b00000011011110000110010001001000;
   assign mem[13916] = 32'b00000001010000100001100110110010;
   assign mem[13917] = 32'b00000001011100010100000100011000;
   assign mem[13918] = 32'b00000000100111001001011111001110;
   assign mem[13919] = 32'b11111101100000111011110000010000;
   assign mem[13920] = 32'b00001000000000011001100010000000;
   assign mem[13921] = 32'b11111011101001001110010101110000;
   assign mem[13922] = 32'b00000101110010001001000000011000;
   assign mem[13923] = 32'b11111111100100000000110000000100;
   assign mem[13924] = 32'b00000010111010011000001011110000;
   assign mem[13925] = 32'b00000010110111110010001111011000;
   assign mem[13926] = 32'b11111110110101010011110100111000;
   assign mem[13927] = 32'b11110111111111111100110111100000;
   assign mem[13928] = 32'b11111001011000010111100111111000;
   assign mem[13929] = 32'b11111001111101111001100001100000;
   assign mem[13930] = 32'b11110001111110101010110011010000;
   assign mem[13931] = 32'b11111110001011000101000110000000;
   assign mem[13932] = 32'b00000010000100111110111110111000;
   assign mem[13933] = 32'b11111110110101100100100100000100;
   assign mem[13934] = 32'b11111101101000001101001110000000;
   assign mem[13935] = 32'b00000000100101001000011110010111;
   assign mem[13936] = 32'b11111001100100011011111011110000;
   assign mem[13937] = 32'b11111111011101101101110011110011;
   assign mem[13938] = 32'b11111100011000111000110111100100;
   assign mem[13939] = 32'b00000101110001001111000001010000;
   assign mem[13940] = 32'b00000101001010101010100011010000;
   assign mem[13941] = 32'b11111111000101001010001100001100;
   assign mem[13942] = 32'b11111101110000111111001011111000;
   assign mem[13943] = 32'b11111100000001111110101110100000;
   assign mem[13944] = 32'b00000110011111100001110011100000;
   assign mem[13945] = 32'b11111011100101010100010110011000;
   assign mem[13946] = 32'b11111100100011010000011010101000;
   assign mem[13947] = 32'b00000101100100010000000111001000;
   assign mem[13948] = 32'b11111100100101100000110000000000;
   assign mem[13949] = 32'b00000011101010110000000111110000;
   assign mem[13950] = 32'b00000011101000101101000111100000;
   assign mem[13951] = 32'b00000100100101011101100111011000;
   assign mem[13952] = 32'b00000011110000101000101001100100;
   assign mem[13953] = 32'b11111111101010000110010000011011;
   assign mem[13954] = 32'b00000010000000101010001001001000;
   assign mem[13955] = 32'b11111110100011011011001000000010;
   assign mem[13956] = 32'b00000010010100111001111000100100;
   assign mem[13957] = 32'b11111010101011100101011101000000;
   assign mem[13958] = 32'b00000010110000100001010101110100;
   assign mem[13959] = 32'b11111010110011101100000100101000;
   assign mem[13960] = 32'b00000100110000110111001011010000;
   assign mem[13961] = 32'b00000011100011101111001010110100;
   assign mem[13962] = 32'b00000011011001010110101110000100;
   assign mem[13963] = 32'b00000001101110000110010101111000;
   assign mem[13964] = 32'b11111110011100000010010101110010;
   assign mem[13965] = 32'b00000011100100101100001100000000;
   assign mem[13966] = 32'b00000010111111111100010011010100;
   assign mem[13967] = 32'b11110100101111011110000100110000;
   assign mem[13968] = 32'b00000010110000101001011110010000;
   assign mem[13969] = 32'b11111010111111100100000110001000;
   assign mem[13970] = 32'b11111111010101001100100011111110;
   assign mem[13971] = 32'b00000101110000110111110000011000;
   assign mem[13972] = 32'b00000000001111010011100111100101;
   assign mem[13973] = 32'b11111111011100101110001001111000;
   assign mem[13974] = 32'b11111011100000001111111000100000;
   assign mem[13975] = 32'b00000011100011111000000011011100;
   assign mem[13976] = 32'b11111100101100000001010001111100;
   assign mem[13977] = 32'b11111110111010111111100001001110;
   assign mem[13978] = 32'b00000010101111011100011111000000;
   assign mem[13979] = 32'b11111110000001010100101101100000;
   assign mem[13980] = 32'b11111111111111111010001100101010;
   assign mem[13981] = 32'b00000000101111111101100111001111;
   assign mem[13982] = 32'b00000110110111000010000111111000;
   assign mem[13983] = 32'b11111110001011001101000000111010;
   assign mem[13984] = 32'b11111010011011010000010011000000;
   assign mem[13985] = 32'b00000100110001000000110100001000;
   assign mem[13986] = 32'b11111111010011110011111110111100;
   assign mem[13987] = 32'b11110110110100110101101101000000;
   assign mem[13988] = 32'b11111110110001100111010111101110;
   assign mem[13989] = 32'b11111101001110110110101111101100;
   assign mem[13990] = 32'b00000100011000100110010110001000;
   assign mem[13991] = 32'b00001101010011100011011011100000;
   assign mem[13992] = 32'b11111100010100111011110110001000;
   assign mem[13993] = 32'b11110101110000001010000110110000;
   assign mem[13994] = 32'b00000010100110111110011001000000;
   assign mem[13995] = 32'b11111000100000111000101100110000;
   assign mem[13996] = 32'b11110110101100001111111011000000;
   assign mem[13997] = 32'b00000110111110110001010110000000;
   assign mem[13998] = 32'b11111110111111111000010001101000;
   assign mem[13999] = 32'b00000110011110101000100001011000;
   assign mem[14000] = 32'b00000100000110001011010111111000;
   assign mem[14001] = 32'b00000000110011110100100010000101;
   assign mem[14002] = 32'b00000011011010110111110111010000;
   assign mem[14003] = 32'b00000100000011100110010100110000;
   assign mem[14004] = 32'b11111001001000011011110001101000;
   assign mem[14005] = 32'b00000100010000110001001010010000;
   assign mem[14006] = 32'b11111111101110101011100101001100;
   assign mem[14007] = 32'b00000101001001111001100011010000;
   assign mem[14008] = 32'b00000010010100110000010111111000;
   assign mem[14009] = 32'b11111001011101111110001011010000;
   assign mem[14010] = 32'b00000001110100110001101000001000;
   assign mem[14011] = 32'b11111011101100100100110010110000;
   assign mem[14012] = 32'b11111101111001011100100001100100;
   assign mem[14013] = 32'b00000000101111100011001110010001;
   assign mem[14014] = 32'b11111100100001010001101110101100;
   assign mem[14015] = 32'b00000010000111100101001101001100;
   assign mem[14016] = 32'b00000011001111000110001011111100;
   assign mem[14017] = 32'b11111110100110011111110011100110;
   assign mem[14018] = 32'b11111110011111010011011100110000;
   assign mem[14019] = 32'b00000000101100010010110101100101;
   assign mem[14020] = 32'b00000000000010010101010011010110;
   assign mem[14021] = 32'b00000101010100110000000111000000;
   assign mem[14022] = 32'b11110111001101011110100100000000;
   assign mem[14023] = 32'b00001010011111010111100011100000;
   assign mem[14024] = 32'b11110010101110101100111110010000;
   assign mem[14025] = 32'b00001000110011001010001100000000;
   assign mem[14026] = 32'b11111000100101111100010001101000;
   assign mem[14027] = 32'b11101111001010011010111101000000;
   assign mem[14028] = 32'b11110001010101010000101101100000;
   assign mem[14029] = 32'b00001000001010011111111101010000;
   assign mem[14030] = 32'b00001001001011000010101011010000;
   assign mem[14031] = 32'b11111001110000001001111000110000;
   assign mem[14032] = 32'b00000101001011100001100101101000;
   assign mem[14033] = 32'b00000010101100000111010000001100;
   assign mem[14034] = 32'b11111000110100011101000100010000;
   assign mem[14035] = 32'b00000100110100001010011111000000;
   assign mem[14036] = 32'b11111110101010010010011010010010;
   assign mem[14037] = 32'b11110100111010110111001100100000;
   assign mem[14038] = 32'b11110011110010110110011001010000;
   assign mem[14039] = 32'b00000010101110010110010011100000;
   assign mem[14040] = 32'b11101000001110111010001111100000;
   assign mem[14041] = 32'b00000100100101001100010101000000;
   assign mem[14042] = 32'b11111110000101010001010110001110;
   assign mem[14043] = 32'b00001010110001101111010110000000;
   assign mem[14044] = 32'b00000010110010001001011111111100;
   assign mem[14045] = 32'b00001111001110100100100110010000;
   assign mem[14046] = 32'b11101101100110111110100000100000;
   assign mem[14047] = 32'b11111111110110101101010100110110;
   assign mem[14048] = 32'b11101010100111010001100001100000;
   assign mem[14049] = 32'b00000101101001101011110011101000;
   assign mem[14050] = 32'b11110011011111111010001101000000;
   assign mem[14051] = 32'b00000001010011010111010000001000;
   assign mem[14052] = 32'b11111110000111010010000111000110;
   assign mem[14053] = 32'b11111000011110110110101101000000;
   assign mem[14054] = 32'b00000101001100111001101011110000;
   assign mem[14055] = 32'b11111111100101100001100101100001;
   assign mem[14056] = 32'b11111000100000010011110011101000;
   assign mem[14057] = 32'b00000111101111001100000001111000;
   assign mem[14058] = 32'b11111010110111110101000000000000;
   assign mem[14059] = 32'b00000110000001001100101011101000;
   assign mem[14060] = 32'b00001000101011000111010110000000;
   assign mem[14061] = 32'b00000010000001101011101000111000;
   assign mem[14062] = 32'b00000101111011000000000011111000;
   assign mem[14063] = 32'b11111111100101100001101111011111;
   assign mem[14064] = 32'b11111011011111000101001010100000;
   assign mem[14065] = 32'b11111110110101101110010011111000;
   assign mem[14066] = 32'b11111110111000100001111011011000;
   assign mem[14067] = 32'b11111101101011000011001001001000;
   assign mem[14068] = 32'b00000110100101001011110111101000;
   assign mem[14069] = 32'b11111011011011110001010000000000;
   assign mem[14070] = 32'b00000011100010110111001101000000;
   assign mem[14071] = 32'b00000101011000011110100011001000;
   assign mem[14072] = 32'b11111111110110000000111000011010;
   assign mem[14073] = 32'b11101111011010100111011111100000;
   assign mem[14074] = 32'b11111110000101101011100110110010;
   assign mem[14075] = 32'b11110100001011010011110111010000;
   assign mem[14076] = 32'b11111001110011111010010000101000;
   assign mem[14077] = 32'b00000000101100100001011011111101;
   assign mem[14078] = 32'b00000100000011111110011101111000;
   assign mem[14079] = 32'b00000000001110010001000010110111;
   assign mem[14080] = 32'b00000110011101011001100110101000;
   assign mem[14081] = 32'b11110101111101111001011111000000;
   assign mem[14082] = 32'b11111011101010010010100001000000;
   assign mem[14083] = 32'b11111010110111001100010001100000;
   assign mem[14084] = 32'b11111110011100001000000100010000;
   assign mem[14085] = 32'b11111011100011011001100100001000;
   assign mem[14086] = 32'b11111110000000011001111001000100;
   assign mem[14087] = 32'b11111111101000111111111010001000;
   assign mem[14088] = 32'b00000010100010111110000111010000;
   assign mem[14089] = 32'b00000110011101010101101100110000;
   assign mem[14090] = 32'b00001111101000101010110111110000;
   assign mem[14091] = 32'b00001100111010001010011010000000;
   assign mem[14092] = 32'b11100010001010110101110100000000;
   assign mem[14093] = 32'b00000001000110100011001010101100;
   assign mem[14094] = 32'b11111011001000001111001100010000;
   assign mem[14095] = 32'b00000010110100111110011101001000;
   assign mem[14096] = 32'b00000000010011011110001101001111;
   assign mem[14097] = 32'b00000100011110101011110001011000;
   assign mem[14098] = 32'b11110011001011111110001010110000;
   assign mem[14099] = 32'b00000100010010100011000101001000;
   assign mem[14100] = 32'b00000111000011000111011111000000;
   assign mem[14101] = 32'b11111010011000111000011010000000;
   assign mem[14102] = 32'b00000110110110010011000011110000;
   assign mem[14103] = 32'b00000100010011001101100011001000;
   assign mem[14104] = 32'b11110100010011101111101110100000;
   assign mem[14105] = 32'b00000001000011101001101101011010;
   assign mem[14106] = 32'b00000111000110001010000110010000;
   assign mem[14107] = 32'b11110100010010000110110011000000;
   assign mem[14108] = 32'b00000011101001111110011110111000;
   assign mem[14109] = 32'b11111110110010001000101011111100;
   assign mem[14110] = 32'b11111101110100001100001101101000;
   assign mem[14111] = 32'b11111110010010111000011100000110;
   assign mem[14112] = 32'b11111100100010110000101011110100;
   assign mem[14113] = 32'b00000000101111111001110010000111;
   assign mem[14114] = 32'b11111101010010010110011000111000;
   assign mem[14115] = 32'b11111111111000110111101001110100;
   assign mem[14116] = 32'b00000011000010100110111000011100;
   assign mem[14117] = 32'b11111010011111100010110001011000;
   assign mem[14118] = 32'b11111111101111011101011110111110;
   assign mem[14119] = 32'b11111110001111010111010110100100;
   assign mem[14120] = 32'b00000000101110001111100111000001;
   assign mem[14121] = 32'b11111010110111111100000100100000;
   assign mem[14122] = 32'b00000111010111011101010011100000;
   assign mem[14123] = 32'b00000000011111100011000101010010;
   assign mem[14124] = 32'b11111011001111111000110110000000;
   assign mem[14125] = 32'b00000010100101111110100011000100;
   assign mem[14126] = 32'b00000011000010100100110001011000;
   assign mem[14127] = 32'b11110111010100010110011000100000;
   assign mem[14128] = 32'b11110111100110100000000111010000;
   assign mem[14129] = 32'b11111111101001110001101101110110;
   assign mem[14130] = 32'b00000010110000010010000111011000;
   assign mem[14131] = 32'b00000000111101010010110100101111;
   assign mem[14132] = 32'b11111011000101001100100100010000;
   assign mem[14133] = 32'b00000000001000100110011011101001;
   assign mem[14134] = 32'b00000100111110111000010110111000;
   assign mem[14135] = 32'b11111110001011010111001010000000;
   assign mem[14136] = 32'b11111101101101001110101111010000;
   assign mem[14137] = 32'b00000101000010101110000010100000;
   assign mem[14138] = 32'b11110111101010011010001100010000;
   assign mem[14139] = 32'b00000010101100111011100100111000;
   assign mem[14140] = 32'b11111000010011010101100001101000;
   assign mem[14141] = 32'b00001010001100111010101110000000;
   assign mem[14142] = 32'b11111100011110011100010010110000;
   assign mem[14143] = 32'b11110001011011000000111101110000;
   assign mem[14144] = 32'b00000100111110110001010000010000;
   assign mem[14145] = 32'b00000111101011111110011011010000;
   assign mem[14146] = 32'b11110011011101000111101010100000;
   assign mem[14147] = 32'b00000100010111111111111101101000;
   assign mem[14148] = 32'b11111101000001110110001010010000;
   assign mem[14149] = 32'b00001001101011101011110101110000;
   assign mem[14150] = 32'b00000111100110110000011111100000;
   assign mem[14151] = 32'b11111100010111110110011001000000;
   assign mem[14152] = 32'b11111110010010101001100101010100;
   assign mem[14153] = 32'b00000011000011001011111010100100;
   assign mem[14154] = 32'b00000001110000110110010110010110;
   assign mem[14155] = 32'b00000100101110001011100100111000;
   assign mem[14156] = 32'b11111110110010000000100000111110;
   assign mem[14157] = 32'b11111110100011011000110110101100;
   assign mem[14158] = 32'b11111001000111100001111101010000;
   assign mem[14159] = 32'b00000010000100111001101010111000;
   assign mem[14160] = 32'b11111110111101100010111000100100;
   assign mem[14161] = 32'b00001101110100011111100111010000;
   assign mem[14162] = 32'b11101110000000101100100000100000;
   assign mem[14163] = 32'b11111111011101111010111001101111;
   assign mem[14164] = 32'b11100110111101001001111101100000;
   assign mem[14165] = 32'b00000100001010000100001011101000;
   assign mem[14166] = 32'b00000011011011110111011110001100;
   assign mem[14167] = 32'b11110111110000011101001011100000;
   assign mem[14168] = 32'b11110111111010011101110101010000;
   assign mem[14169] = 32'b00000101000000111000010100001000;
   assign mem[14170] = 32'b11100110000110100110100110100000;
   assign mem[14171] = 32'b00000101011100001100101001001000;
   assign mem[14172] = 32'b00000000001011000101111010101001;
   assign mem[14173] = 32'b11110111000110100100001100000000;
   assign mem[14174] = 32'b00000011001110011000110001101000;
   assign mem[14175] = 32'b11111001101011011000100111100000;
   assign mem[14176] = 32'b11100100111000101011000010000000;
   assign mem[14177] = 32'b00000110010110110011010000111000;
   assign mem[14178] = 32'b11111010011001001010100101110000;
   assign mem[14179] = 32'b00000111000110101110111011001000;
   assign mem[14180] = 32'b00000010111000000010010010101000;
   assign mem[14181] = 32'b00001000011110010110111100000000;
   assign mem[14182] = 32'b11111100010011011000101110111000;
   assign mem[14183] = 32'b00000000010011101000011001010010;
   assign mem[14184] = 32'b11111100000000000101011000100100;
   assign mem[14185] = 32'b00000001011000010100101011110000;
   assign mem[14186] = 32'b00000010001000100111010110101000;
   assign mem[14187] = 32'b11110111101110111010100011100000;
   assign mem[14188] = 32'b00000001001101000011001011110010;
   assign mem[14189] = 32'b00000011110000000001010100101000;
   assign mem[14190] = 32'b00000110111100101011111001111000;
   assign mem[14191] = 32'b11111010000010000011100110001000;
   assign mem[14192] = 32'b11111111101011101101000011100011;
   assign mem[14193] = 32'b11111011001111101001011011011000;
   assign mem[14194] = 32'b11111010000000000101100000100000;
   assign mem[14195] = 32'b00000001000110001010101101101010;
   assign mem[14196] = 32'b00000011101010101001111100110100;
   assign mem[14197] = 32'b11111010101111001010010100010000;
   assign mem[14198] = 32'b00000010101101111010111011011000;
   assign mem[14199] = 32'b00000000110110001000111011111111;
   assign mem[14200] = 32'b00000001011110001110011110111100;
   assign mem[14201] = 32'b00000100100010010001101000001000;
   assign mem[14202] = 32'b00000100110000111111001011101000;
   assign mem[14203] = 32'b11110111000101111110110000110000;
   assign mem[14204] = 32'b00000110011010001001110100110000;
   assign mem[14205] = 32'b11111110110111001111010100110100;
   assign mem[14206] = 32'b11111001001101100111001001010000;
   assign mem[14207] = 32'b11111001110100100100111110010000;
   assign mem[14208] = 32'b11111111000010101101010010010101;
   assign mem[14209] = 32'b00000011010100100011100010111100;
   assign mem[14210] = 32'b00000101010010100001111110101000;
   assign mem[14211] = 32'b11111001100001001011000010010000;
   assign mem[14212] = 32'b00000000111001110001010100100010;
   assign mem[14213] = 32'b00000000010010110001101010011111;
   assign mem[14214] = 32'b11111011001101010000100000111000;
   assign mem[14215] = 32'b00000110001110010010100100101000;
   assign mem[14216] = 32'b00000010101001110100101001010100;
   assign mem[14217] = 32'b11111000101101010110011101100000;
   assign mem[14218] = 32'b00000001011010010100100100010110;
   assign mem[14219] = 32'b11111110110110111001010001110100;
   assign mem[14220] = 32'b00000011100110111000111001111000;
   assign mem[14221] = 32'b11111101101000110111101101010100;
   assign mem[14222] = 32'b00001000010111010010011000110000;
   assign mem[14223] = 32'b11111101111001010100100010110100;
   assign mem[14224] = 32'b11111011001111100000101001100000;
   assign mem[14225] = 32'b11111111001010011010000111000001;
   assign mem[14226] = 32'b00000010101010111111011101001100;
   assign mem[14227] = 32'b11111100001000100011110001011000;
   assign mem[14228] = 32'b00000111000000011001001110101000;
   assign mem[14229] = 32'b11111000010110100000100110000000;
   assign mem[14230] = 32'b11110110101010010100010000110000;
   assign mem[14231] = 32'b00000101001011001000010110011000;
   assign mem[14232] = 32'b11110111000110101011011000110000;
   assign mem[14233] = 32'b00000100111110011110111101011000;
   assign mem[14234] = 32'b00000011011110101010011000010000;
   assign mem[14235] = 32'b00000010110011111101000010011000;
   assign mem[14236] = 32'b11101111101100000101010101100000;
   assign mem[14237] = 32'b00000101000001100101010111000000;
   assign mem[14238] = 32'b11111001000111101110011001001000;
   assign mem[14239] = 32'b00000100010100000111001111011000;
   assign mem[14240] = 32'b00000101001001011001011011101000;
   assign mem[14241] = 32'b00000000110011001101010010011101;
   assign mem[14242] = 32'b00000101001111011110011101100000;
   assign mem[14243] = 32'b00000000110010010010110001001100;
   assign mem[14244] = 32'b11111011111001110011110111011000;
   assign mem[14245] = 32'b00000001111010011001100000101100;
   assign mem[14246] = 32'b00000011110111010011010110000100;
   assign mem[14247] = 32'b11110100001100010001011001000000;
   assign mem[14248] = 32'b00000010010111011101010101001100;
   assign mem[14249] = 32'b11111100011001001000000000010100;
   assign mem[14250] = 32'b11111100000110001010100101100100;
   assign mem[14251] = 32'b00001001110000110110100011000000;
   assign mem[14252] = 32'b00000010101101010000101000010100;
   assign mem[14253] = 32'b11111000010100011000111001101000;
   assign mem[14254] = 32'b00000000100011110101111101010111;
   assign mem[14255] = 32'b11111111100000110011101000001100;
   assign mem[14256] = 32'b00000101100001100111100010100000;
   assign mem[14257] = 32'b11111100101011000100000110111000;
   assign mem[14258] = 32'b00000001001011011110111111101110;
   assign mem[14259] = 32'b11111111001000111111110101000100;
   assign mem[14260] = 32'b00000010111100111111001000011100;
   assign mem[14261] = 32'b00001100111001001011011000100000;
   assign mem[14262] = 32'b00000101100110001111010000010000;
   assign mem[14263] = 32'b11111100110011110100110101101000;
   assign mem[14264] = 32'b11111010011011100011111010100000;
   assign mem[14265] = 32'b11111110111100001000000110000000;
   assign mem[14266] = 32'b11111101011010111100001000011100;
   assign mem[14267] = 32'b11110000000011001000110011000000;
   assign mem[14268] = 32'b11111100101100111101000101101000;
   assign mem[14269] = 32'b11111011101101010000001111011000;
   assign mem[14270] = 32'b11110110111000111010011110010000;
   assign mem[14271] = 32'b11110010100000011001011111010000;
   assign mem[14272] = 32'b00000111000001001011111110101000;
   assign mem[14273] = 32'b00001001110001010110110010010000;
   assign mem[14274] = 32'b11110111110110110010100000010000;
   assign mem[14275] = 32'b00000000011010011001001100000111;
   assign mem[14276] = 32'b11110101010111101010010001000000;
   assign mem[14277] = 32'b11101110001000010000101000100000;
   assign mem[14278] = 32'b00000010001000010010111100101000;
   assign mem[14279] = 32'b00000000100001110001111101111110;
   assign mem[14280] = 32'b11101100000011101111000000100000;
   assign mem[14281] = 32'b00000110101101101011010111101000;
   assign mem[14282] = 32'b11111100000011011100010011110000;
   assign mem[14283] = 32'b11110100010110010010000100010000;
   assign mem[14284] = 32'b00000110010001101110111010100000;
   assign mem[14285] = 32'b11110001110000010011011111100000;
   assign mem[14286] = 32'b11110010100111001001010000110000;
   assign mem[14287] = 32'b00000100010000101100000111010000;
   assign mem[14288] = 32'b00000010110100011110000000110100;
   assign mem[14289] = 32'b00000110000101000101101101011000;
   assign mem[14290] = 32'b00000000011110100010010000110011;
   assign mem[14291] = 32'b11111110010111111111100101001110;
   assign mem[14292] = 32'b00000001111110010110100110111010;
   assign mem[14293] = 32'b00000101011000010000010001101000;
   assign mem[14294] = 32'b11111000100100110110101111011000;
   assign mem[14295] = 32'b00000100101101000011100101010000;
   assign mem[14296] = 32'b11111110111110010000110101110000;
   assign mem[14297] = 32'b11100011000111101111110111000000;
   assign mem[14298] = 32'b00000001100100001011100111011010;
   assign mem[14299] = 32'b11111100111011110111100000101100;
   assign mem[14300] = 32'b00000111000011100000001110010000;
   assign mem[14301] = 32'b11110110010011000101000100110000;
   assign mem[14302] = 32'b11111001010110100000001101001000;
   assign mem[14303] = 32'b00001000001010010011111111000000;
   assign mem[14304] = 32'b00000100010011100110001111010000;
   assign mem[14305] = 32'b00000011001110010011111000000100;
   assign mem[14306] = 32'b11111100010100001000001001010000;
   assign mem[14307] = 32'b00000011110111010010100110000100;
   assign mem[14308] = 32'b11111100010110111011101111100000;
   assign mem[14309] = 32'b00000101011010001011001101011000;
   assign mem[14310] = 32'b00000110101010111110001100001000;
   assign mem[14311] = 32'b00000001010001000000101110000000;
   assign mem[14312] = 32'b00000000111001010111010111000110;
   assign mem[14313] = 32'b11111111001100010101101010001101;
   assign mem[14314] = 32'b11111000000111000100000111100000;
   assign mem[14315] = 32'b11111100001101101010001110111100;
   assign mem[14316] = 32'b00000101100111110100111011101000;
   assign mem[14317] = 32'b11111101111000101010111010000100;
   assign mem[14318] = 32'b00000001101111001111000010110000;
   assign mem[14319] = 32'b11111100110110101101111111011000;
   assign mem[14320] = 32'b00001001110101100100011000100000;
   assign mem[14321] = 32'b00000000001011011111010100111111;
   assign mem[14322] = 32'b11111011100010000000000111100000;
   assign mem[14323] = 32'b11111010100111001010011101111000;
   assign mem[14324] = 32'b11111110111000100110010100011100;
   assign mem[14325] = 32'b11111111000111100110011001001010;
   assign mem[14326] = 32'b00000100000000110011111000110000;
   assign mem[14327] = 32'b11111101111011101110001101100000;
   assign mem[14328] = 32'b00000011001011101111110100100000;
   assign mem[14329] = 32'b11111011101110001011101101110000;
   assign mem[14330] = 32'b11110001101010001111100101010000;
   assign mem[14331] = 32'b00001000101110101100000110000000;
   assign mem[14332] = 32'b11110110100110000100000100110000;
   assign mem[14333] = 32'b11110000000001000011000101110000;
   assign mem[14334] = 32'b00000101101110011010110011110000;
   assign mem[14335] = 32'b00001000010011011100000111100000;
   assign mem[14336] = 32'b11101111111000011001110101100000;
   assign mem[14337] = 32'b00000111100000101101101100010000;
   assign mem[14338] = 32'b11111011001001010111010011010000;
   assign mem[14339] = 32'b00000101111001001000000100111000;
   assign mem[14340] = 32'b00000101101101100101110111000000;
   assign mem[14341] = 32'b00000011001010001101100010000100;
   assign mem[14342] = 32'b11111101010111001110010100110100;
   assign mem[14343] = 32'b11100111110011011100010110000000;
   assign mem[14344] = 32'b00000000100110001010001101101100;
   assign mem[14345] = 32'b11111000001010100000101010011000;
   assign mem[14346] = 32'b00000001001101001111101010100010;
   assign mem[14347] = 32'b00000010110111010110010001100000;
   assign mem[14348] = 32'b00000101101010000111101010100000;
   assign mem[14349] = 32'b11111111010010111010100111011000;
   assign mem[14350] = 32'b11111001101100010100001111111000;
   assign mem[14351] = 32'b00001111110111100000111100110000;
   assign mem[14352] = 32'b00000111110001111010001011100000;
   assign mem[14353] = 32'b00001001011111010111110110110000;
   assign mem[14354] = 32'b11110100101001110011110111110000;
   assign mem[14355] = 32'b00000111000111011001101101110000;
   assign mem[14356] = 32'b11101101101101000001010001000000;
   assign mem[14357] = 32'b00000011010001111011011111000100;
   assign mem[14358] = 32'b11110110001001111100000110100000;
   assign mem[14359] = 32'b11111101011000111110110101000000;
   assign mem[14360] = 32'b00000100101101110011101011001000;
   assign mem[14361] = 32'b11111000100111110110001011100000;
   assign mem[14362] = 32'b00000010000010011011100001011000;
   assign mem[14363] = 32'b00000001110100011111111011000010;
   assign mem[14364] = 32'b11111011010110001111111110100000;
   assign mem[14365] = 32'b00000000000111110010001111011010;
   assign mem[14366] = 32'b00000010111100001101111011101100;
   assign mem[14367] = 32'b11111001010011001000010100100000;
   assign mem[14368] = 32'b00000101010010100001101111001000;
   assign mem[14369] = 32'b11111100001010010101111101001100;
   assign mem[14370] = 32'b11111101111000011011100000111000;
   assign mem[14371] = 32'b00001000010111100111110101110000;
   assign mem[14372] = 32'b11110110001010000010111111000000;
   assign mem[14373] = 32'b00000000011110100111010001100001;
   assign mem[14374] = 32'b11110001101101001010001100100000;
   assign mem[14375] = 32'b00000011100001000111001100011000;
   assign mem[14376] = 32'b11111100110010100011000111011100;
   assign mem[14377] = 32'b11111100010101100101011101001100;
   assign mem[14378] = 32'b11111010011111011011111010111000;
   assign mem[14379] = 32'b11111111110010011010110011010011;
   assign mem[14380] = 32'b11110100101101100101001111000000;
   assign mem[14381] = 32'b00001010001010110011011100010000;
   assign mem[14382] = 32'b11110110001110000010000000100000;
   assign mem[14383] = 32'b11111101101001110110110101000100;
   assign mem[14384] = 32'b00000101000011010000011101110000;
   assign mem[14385] = 32'b11111100010110101011000001001000;
   assign mem[14386] = 32'b11110110001000100110000101000000;
   assign mem[14387] = 32'b00000100100101011001110011111000;
   assign mem[14388] = 32'b00000000001111010111111010001101;
   assign mem[14389] = 32'b00000111110111100100110001011000;
   assign mem[14390] = 32'b00000001100010011000011111001010;
   assign mem[14391] = 32'b11111111100111001010101101111101;
   assign mem[14392] = 32'b11111100100000000001001111010000;
   assign mem[14393] = 32'b00000000101010010011001110100100;
   assign mem[14394] = 32'b11111110100010011011111110111000;
   assign mem[14395] = 32'b11111101110100001101100111001000;
   assign mem[14396] = 32'b00000000001011000111111111011001;
   assign mem[14397] = 32'b11111011101110110010001101001000;
   assign mem[14398] = 32'b11111111101000111010010100010110;
   assign mem[14399] = 32'b00000001100001100110001110011110;
   assign mem[14400] = 32'b00000100110111101111111010100000;
   assign mem[14401] = 32'b00000001110110000011011010011100;
   assign mem[14402] = 32'b00000010001110111011100011111000;
   assign mem[14403] = 32'b00000111001000110101101011011000;
   assign mem[14404] = 32'b11111101100101001001111010010100;
   assign mem[14405] = 32'b00000011010111000010101010111000;
   assign mem[14406] = 32'b11111010101101111001001001100000;
   assign mem[14407] = 32'b11111011000001110011101110110000;
   assign mem[14408] = 32'b11110010111110000011100101110000;
   assign mem[14409] = 32'b11111111110000101111011111110101;
   assign mem[14410] = 32'b11111100100011010100000110111000;
   assign mem[14411] = 32'b00000010010000001010010111111000;
   assign mem[14412] = 32'b11111000110110001011011111111000;
   assign mem[14413] = 32'b00000001001011011001110100100110;
   assign mem[14414] = 32'b00000100000000000110000111011000;
   assign mem[14415] = 32'b11111010100010010111000010101000;
   assign mem[14416] = 32'b11110110101101001011010000110000;
   assign mem[14417] = 32'b00000101101000000010111011010000;
   assign mem[14418] = 32'b11110110111000010101100011100000;
   assign mem[14419] = 32'b00000100100000110110100110001000;
   assign mem[14420] = 32'b00000001010100101001100010001100;
   assign mem[14421] = 32'b00000011010110101001001010110000;
   assign mem[14422] = 32'b00000000111100000010101101000100;
   assign mem[14423] = 32'b11111101111011000101101101100000;
   assign mem[14424] = 32'b11111000010000101111101011000000;
   assign mem[14425] = 32'b00000000001101111001000100010110;
   assign mem[14426] = 32'b00000011010001000001111100000000;
   assign mem[14427] = 32'b11111101011110010010110010010000;
   assign mem[14428] = 32'b11111111100001000101010010101101;
   assign mem[14429] = 32'b11111100001011001010110001010000;
   assign mem[14430] = 32'b11111100001011101010110111100000;
   assign mem[14431] = 32'b00001000100001011000001100000000;
   assign mem[14432] = 32'b11111010000000101101100110011000;
   assign mem[14433] = 32'b11110111000110000010110111100000;
   assign mem[14434] = 32'b11111110000110110101001110001010;
   assign mem[14435] = 32'b00001100100111010101011010110000;
   assign mem[14436] = 32'b11110110101011000001011101010000;
   assign mem[14437] = 32'b00000011101101101100110110100100;
   assign mem[14438] = 32'b11111111100101001110010001011110;
   assign mem[14439] = 32'b00000011000111100010000001101100;
   assign mem[14440] = 32'b00001000100000010001110110010000;
   assign mem[14441] = 32'b11110111010101101101101000010000;
   assign mem[14442] = 32'b00000011010001010101111000010100;
   assign mem[14443] = 32'b00000100011100111000001000100000;
   assign mem[14444] = 32'b11111000110011001110001010011000;
   assign mem[14445] = 32'b00000011011011001101010110000100;
   assign mem[14446] = 32'b00000100110101011011001001000000;
   assign mem[14447] = 32'b11101011011110111000101100000000;
   assign mem[14448] = 32'b11111101100010101100000001010000;
   assign mem[14449] = 32'b11111111001000110001111111010001;
   assign mem[14450] = 32'b00000001011111110001110010000100;
   assign mem[14451] = 32'b00001000010010011001111101100000;
   assign mem[14452] = 32'b11111111001000101100101110110011;
   assign mem[14453] = 32'b11111111110100101010101001100100;
   assign mem[14454] = 32'b11110101100001001101110111000000;
   assign mem[14455] = 32'b00000001100110111010111111010010;
   assign mem[14456] = 32'b00000000010011111101011001110101;
   assign mem[14457] = 32'b11110111110110110101011000010000;
   assign mem[14458] = 32'b00000111010001110101010010001000;
   assign mem[14459] = 32'b00000001001011100011111110110000;
   assign mem[14460] = 32'b00001000001011010001001010100000;
   assign mem[14461] = 32'b00000000100101010011010110110110;
   assign mem[14462] = 32'b00000111010001000101011110110000;
   assign mem[14463] = 32'b11111111100010110100001011110010;
   assign mem[14464] = 32'b11111000111110111000001000111000;
   assign mem[14465] = 32'b11111111001101010100111110000001;
   assign mem[14466] = 32'b00000101001010101100100011000000;
   assign mem[14467] = 32'b11111000010110001101100110011000;
   assign mem[14468] = 32'b00000010000110010101110100101000;
   assign mem[14469] = 32'b11110011001101011000010001010000;
   assign mem[14470] = 32'b00000010001011000010110011101100;
   assign mem[14471] = 32'b11110100110110011111011110110000;
   assign mem[14472] = 32'b00000011001101100100001110101100;
   assign mem[14473] = 32'b00001100111000101101111001000000;
   assign mem[14474] = 32'b11110111111110110111000011100000;
   assign mem[14475] = 32'b00001000101010001011100010100000;
   assign mem[14476] = 32'b11111011001010101001000011110000;
   assign mem[14477] = 32'b11110111100001100101001001110000;
   assign mem[14478] = 32'b11101111011010111010010100000000;
   assign mem[14479] = 32'b11111111101001111011101111100111;
   assign mem[14480] = 32'b00000101101011010000111001101000;
   assign mem[14481] = 32'b00000001101010010111010100111100;
   assign mem[14482] = 32'b00000111000011100010101010110000;
   assign mem[14483] = 32'b11111111001010011101101110000001;
   assign mem[14484] = 32'b11110110000111100100110111010000;
   assign mem[14485] = 32'b11111100101010101000000011011100;
   assign mem[14486] = 32'b00000111101010001111111100011000;
   assign mem[14487] = 32'b11110111100110001001111000000000;
   assign mem[14488] = 32'b11111110101011110000100001001100;
   assign mem[14489] = 32'b11111011110100001010111111101000;
   assign mem[14490] = 32'b00000010100110000011101000111000;
   assign mem[14491] = 32'b11111111101010000100001000111101;
   assign mem[14492] = 32'b00000000101011100000000000100111;
   assign mem[14493] = 32'b11111101101010001100101111011100;
   assign mem[14494] = 32'b11111111010001001110011110010011;
   assign mem[14495] = 32'b00000010110001110110100111110100;
   assign mem[14496] = 32'b00000100001110110101010010101000;
   assign mem[14497] = 32'b11110111111001100100010100110000;
   assign mem[14498] = 32'b11111101111110010100111100110100;
   assign mem[14499] = 32'b11111111100100111101111000110010;
   assign mem[14500] = 32'b00000010011010000101111101101000;
   assign mem[14501] = 32'b00000001010111000011110111000110;
   assign mem[14502] = 32'b00000100100100101011011001010000;
   assign mem[14503] = 32'b00000001100101011100110000111100;
   assign mem[14504] = 32'b11111011010001001110111111011000;
   assign mem[14505] = 32'b11111101110110101000111100101100;
   assign mem[14506] = 32'b00000010111001001110011010011000;
   assign mem[14507] = 32'b11111000001000001001011010110000;
   assign mem[14508] = 32'b00000000010100001001101011110001;
   assign mem[14509] = 32'b11111001010011111001000111111000;
   assign mem[14510] = 32'b00010001110100001010001001000000;
   assign mem[14511] = 32'b00000101111100110101000100010000;
   assign mem[14512] = 32'b00000000001000010110000011001110;
   assign mem[14513] = 32'b11111100110000110010001111111100;
   assign mem[14514] = 32'b11110111010101111101110110010000;
   assign mem[14515] = 32'b11111111100110101001010110000001;
   assign mem[14516] = 32'b00000100111010111010011001101000;
   assign mem[14517] = 32'b00000000111101111110101101110001;
   assign mem[14518] = 32'b00000001100101001111110000101110;
   assign mem[14519] = 32'b11110001110011000110101001100000;
   assign mem[14520] = 32'b00001001010001111100111110110000;
   assign mem[14521] = 32'b00000100100000111110111011111000;
   assign mem[14522] = 32'b00000110001100100010011010100000;
   assign mem[14523] = 32'b11111110000111001011100001000100;
   assign mem[14524] = 32'b11110100011011010100011001010000;
   assign mem[14525] = 32'b11111101011000010110011110000000;
   assign mem[14526] = 32'b00000110010010100001011100111000;
   assign mem[14527] = 32'b11111101101110011100011100100100;
   assign mem[14528] = 32'b00000110000010101111000110110000;
   assign mem[14529] = 32'b11101101111010000100111001000000;
   assign mem[14530] = 32'b00000001110100011000111110011010;
   assign mem[14531] = 32'b11111010100001101100010100010000;
   assign mem[14532] = 32'b11111010101100111100111000010000;
   assign mem[14533] = 32'b00000111001001010010101000110000;
   assign mem[14534] = 32'b00000011100111001000011100001100;
   assign mem[14535] = 32'b00001000011101110111101000010000;
   assign mem[14536] = 32'b00000101000010010100011010110000;
   assign mem[14537] = 32'b00000001101101001010101010010010;
   assign mem[14538] = 32'b11110101111100101011010110110000;
   assign mem[14539] = 32'b11111000100100110101100110100000;
   assign mem[14540] = 32'b11110100111100011100010100110000;
   assign mem[14541] = 32'b00001011011101101000101100000000;
   assign mem[14542] = 32'b11110011110101111001110101100000;
   assign mem[14543] = 32'b11110101110100101000000001010000;
   assign mem[14544] = 32'b00000111111011000011100001111000;
   assign mem[14545] = 32'b11110111111100111100000011110000;
   assign mem[14546] = 32'b11110111101010101010000110000000;
   assign mem[14547] = 32'b00001100101100111101101100110000;
   assign mem[14548] = 32'b11110100010101111111100110010000;
   assign mem[14549] = 32'b00001010110111011011010110010000;
   assign mem[14550] = 32'b00000001000001101110101000001100;
   assign mem[14551] = 32'b11111101101100010011001111110000;
   assign mem[14552] = 32'b11111111110101100100111011100010;
   assign mem[14553] = 32'b11111101101110101000111100010000;
   assign mem[14554] = 32'b00000011101000100000010010110100;
   assign mem[14555] = 32'b11111101111000101000100101110000;
   assign mem[14556] = 32'b11111100001100101010010000111000;
   assign mem[14557] = 32'b00000011100010010100011111000000;
   assign mem[14558] = 32'b00000010111001001000110100001000;
   assign mem[14559] = 32'b11111100100000111110100011111100;
   assign mem[14560] = 32'b00000000110110100110001110100000;
   assign mem[14561] = 32'b00000000011011000001101010100100;
   assign mem[14562] = 32'b00000110000001101101011000100000;
   assign mem[14563] = 32'b00000001000010111010011000100100;
   assign mem[14564] = 32'b11111101000000001101010001000100;
   assign mem[14565] = 32'b00000110000001010110001110101000;
   assign mem[14566] = 32'b00000010001010000001101011000000;
   assign mem[14567] = 32'b11111011101100011110100011101000;
   assign mem[14568] = 32'b11111110111110100000001001111000;
   assign mem[14569] = 32'b11110101100010110111001001000000;
   assign mem[14570] = 32'b11111111011101110000111001000111;
   assign mem[14571] = 32'b00000001000011101110011100010110;
   assign mem[14572] = 32'b00000010001000111100101101010100;
   assign mem[14573] = 32'b00000010111000101111011011101000;
   assign mem[14574] = 32'b11111100011000000000100100001100;
   assign mem[14575] = 32'b00000010111000000011010001110100;
   assign mem[14576] = 32'b11111011100011011110111100100000;
   assign mem[14577] = 32'b11111111010011000000111001100111;
   assign mem[14578] = 32'b11111000001110100000111110111000;
   assign mem[14579] = 32'b00000000000010110000101001001101;
   assign mem[14580] = 32'b00000010010111111011010100000100;
   assign mem[14581] = 32'b11101011100111001100110011000000;
   assign mem[14582] = 32'b00000001011111101110001010100100;
   assign mem[14583] = 32'b00001000001010111000101000100000;
   assign mem[14584] = 32'b11111101101001100110001000011100;
   assign mem[14585] = 32'b00000110001111011011100110100000;
   assign mem[14586] = 32'b11111111000001111110110100100110;
   assign mem[14587] = 32'b11111101001100011011110010110000;
   assign mem[14588] = 32'b00000111001100100111010000101000;
   assign mem[14589] = 32'b11111101001101010100001110010000;
   assign mem[14590] = 32'b11011111011001101010100111000000;
   assign mem[14591] = 32'b00000111111001110001010011001000;
   assign mem[14592] = 32'b11111001001110001100011010011000;
   assign mem[14593] = 32'b11110110011110000001000010110000;
   assign mem[14594] = 32'b00000111010110100000101110000000;
   assign mem[14595] = 32'b11110101011001011111110100010000;
   assign mem[14596] = 32'b11110110001000010111111000010000;
   assign mem[14597] = 32'b00000110011010110101110011011000;
   assign mem[14598] = 32'b11111100000111101011110011001100;
   assign mem[14599] = 32'b00001000100001110100110110100000;
   assign mem[14600] = 32'b11111111111011110000110001100001;
   assign mem[14601] = 32'b00000000101110010000010000001011;
   assign mem[14602] = 32'b11111100101101000111001011011000;
   assign mem[14603] = 32'b11111101100111100111010010011100;
   assign mem[14604] = 32'b11111000110111010011001100100000;
   assign mem[14605] = 32'b11111111110110111111110110010011;
   assign mem[14606] = 32'b00000001101110110110100010001110;
   assign mem[14607] = 32'b11111001001110111010010011011000;
   assign mem[14608] = 32'b00000001101010010011111011111100;
   assign mem[14609] = 32'b11111011101100001101010110111000;
   assign mem[14610] = 32'b11111110100111100011000111111000;
   assign mem[14611] = 32'b00000101000101010111110100010000;
   assign mem[14612] = 32'b00000001100000010000101111111100;
   assign mem[14613] = 32'b00000001000101011110110101101100;
   assign mem[14614] = 32'b11111000111100101010011100100000;
   assign mem[14615] = 32'b11111111110100111100000100100001;
   assign mem[14616] = 32'b00000010101110100000100100000100;
   assign mem[14617] = 32'b11110011010100111110010111000000;
   assign mem[14618] = 32'b00000000000010110111100010000101;
   assign mem[14619] = 32'b11111101100100000100011111000100;
   assign mem[14620] = 32'b00000011010011101110000010011000;
   assign mem[14621] = 32'b00000010010011011011101011010100;
   assign mem[14622] = 32'b11111101100110010101110100001100;
   assign mem[14623] = 32'b00000000101001011100101001101111;
   assign mem[14624] = 32'b11111011110100000101011101111000;
   assign mem[14625] = 32'b00000001011111110110000010011100;
   assign mem[14626] = 32'b00000010000001001000111001010000;
   assign mem[14627] = 32'b11111011000110000001101010000000;
   assign mem[14628] = 32'b11111100100100001100000101011000;
   assign mem[14629] = 32'b11111010101110100010100000110000;
   assign mem[14630] = 32'b11111010110010100110011011111000;
   assign mem[14631] = 32'b00000010100011010000001011111100;
   assign mem[14632] = 32'b11110011110000101100111001100000;
   assign mem[14633] = 32'b11101100111010011111000000000000;
   assign mem[14634] = 32'b00000100010100000010001100111000;
   assign mem[14635] = 32'b00000000010111010000011001010011;
   assign mem[14636] = 32'b11110000010101000011111010000000;
   assign mem[14637] = 32'b00000110100101001000010110001000;
   assign mem[14638] = 32'b00000000100011011001010000110101;
   assign mem[14639] = 32'b00000110000110110110010011000000;
   assign mem[14640] = 32'b11111001101111000010001011010000;
   assign mem[14641] = 32'b00000100011110101000111011010000;
   assign mem[14642] = 32'b11110110111100101001011000010000;
   assign mem[14643] = 32'b00000001111110011110111111001000;
   assign mem[14644] = 32'b11111001000010001000011100011000;
   assign mem[14645] = 32'b00001111000001011011000001110000;
   assign mem[14646] = 32'b00000000101001010000000010100000;
   assign mem[14647] = 32'b11111011011101101111100001000000;
   assign mem[14648] = 32'b00000101000010011111000100011000;
   assign mem[14649] = 32'b11110110111010001011111110000000;
   assign mem[14650] = 32'b00000010110010111101000001011000;
   assign mem[14651] = 32'b11111001111110111111000101011000;
   assign mem[14652] = 32'b11111111000110011111101111101011;
   assign mem[14653] = 32'b11111101100111101001111111111000;
   assign mem[14654] = 32'b00000010101001100100100110110100;
   assign mem[14655] = 32'b00000011001000001100111111010000;
   assign mem[14656] = 32'b00000011010111010111100111000000;
   assign mem[14657] = 32'b11111010111010100110101001100000;
   assign mem[14658] = 32'b11111110011111011001010110000110;
   assign mem[14659] = 32'b11111111101010001100011010100001;
   assign mem[14660] = 32'b00001011100100101110000011000000;
   assign mem[14661] = 32'b11110110100010001101111011110000;
   assign mem[14662] = 32'b11110111100100111000000011010000;
   assign mem[14663] = 32'b00000110111110011100001001100000;
   assign mem[14664] = 32'b11101100110010011011000000100000;
   assign mem[14665] = 32'b00001010010010001010010111010000;
   assign mem[14666] = 32'b11111011101101000000100001100000;
   assign mem[14667] = 32'b11110001001011111010011010000000;
   assign mem[14668] = 32'b11110101101100000010101111110000;
   assign mem[14669] = 32'b00000100110011100101011100001000;
   assign mem[14670] = 32'b00000100110011100111110100000000;
   assign mem[14671] = 32'b00000010010110111001101110100000;
   assign mem[14672] = 32'b11111001101001101011010101111000;
   assign mem[14673] = 32'b00001010001001101010101111000000;
   assign mem[14674] = 32'b11101100001001110111010100000000;
   assign mem[14675] = 32'b00000111100101111011010101100000;
   assign mem[14676] = 32'b00000001100000011111100101010110;
   assign mem[14677] = 32'b11110101111000101111111111100000;
   assign mem[14678] = 32'b11111111100111010100000010010111;
   assign mem[14679] = 32'b11110101111001110100000001000000;
   assign mem[14680] = 32'b11110100100100100111100010010000;
   assign mem[14681] = 32'b00001010110011001001001110110000;
   assign mem[14682] = 32'b00000001011000111000110001000100;
   assign mem[14683] = 32'b00010001000011011001101110000000;
   assign mem[14684] = 32'b11110100110111000110001001110000;
   assign mem[14685] = 32'b00000111101010000110101010001000;
   assign mem[14686] = 32'b11100111111101101000101100000000;
   assign mem[14687] = 32'b11111010000000110111010101100000;
   assign mem[14688] = 32'b11101110100010111100000100000000;
   assign mem[14689] = 32'b00000100101101011111111011100000;
   assign mem[14690] = 32'b11111100111000000010111001101100;
   assign mem[14691] = 32'b00000010001010011001001101100100;
   assign mem[14692] = 32'b00000110010011101010000110101000;
   assign mem[14693] = 32'b00000010011001011100011110111100;
   assign mem[14694] = 32'b11111111100100101000000010101000;
   assign mem[14695] = 32'b11111110110101110100101111001010;
   assign mem[14696] = 32'b11111101011000001110010110010000;
   assign mem[14697] = 32'b00000000101010101101000010111110;
   assign mem[14698] = 32'b11110110011011010001111000110000;
   assign mem[14699] = 32'b00000001110000100110010001100000;
   assign mem[14700] = 32'b11111100010110000100111100110100;
   assign mem[14701] = 32'b00000100000001001010011100101000;
   assign mem[14702] = 32'b00000001000111011001100101000000;
   assign mem[14703] = 32'b11110010110111011101001111000000;
   assign mem[14704] = 32'b00000000001010011010011100101001;
   assign mem[14705] = 32'b11101110010011100000010101000000;
   assign mem[14706] = 32'b11110000110010001001011000100000;
   assign mem[14707] = 32'b00000000011010010000000011001110;
   assign mem[14708] = 32'b11111111000111100101101110110000;
   assign mem[14709] = 32'b00000001010110111100010110111000;
   assign mem[14710] = 32'b11111010101001100111001110001000;
   assign mem[14711] = 32'b11111110001001111010001011110000;
   assign mem[14712] = 32'b11111101110000111110010110001000;
   assign mem[14713] = 32'b11111100100111010011011011111000;
   assign mem[14714] = 32'b00000010001011000001110001111100;
   assign mem[14715] = 32'b11111100011010001111111111110000;
   assign mem[14716] = 32'b11101011101101000010001000000000;
   assign mem[14717] = 32'b00000010110000110101101111011000;
   assign mem[14718] = 32'b11111011100010101101001011010000;
   assign mem[14719] = 32'b00000101100010111010000100100000;
   assign mem[14720] = 32'b00000001100010110011010011111010;
   assign mem[14721] = 32'b11101000010100011001000111100000;
   assign mem[14722] = 32'b00001011001010101000100111010000;
   assign mem[14723] = 32'b00000100000101111010001110000000;
   assign mem[14724] = 32'b11111100111011011010011110101100;
   assign mem[14725] = 32'b11111100110010001000011010111100;
   assign mem[14726] = 32'b00001000010100110000101111000000;
   assign mem[14727] = 32'b11111000110110001101111011111000;
   assign mem[14728] = 32'b00000011000100011011000110010100;
   assign mem[14729] = 32'b11111101011000010000011101111100;
   assign mem[14730] = 32'b11011111010100101110110101000000;
   assign mem[14731] = 32'b00000111010000101000011101111000;
   assign mem[14732] = 32'b11110010010100101001110100000000;
   assign mem[14733] = 32'b00000111011001110111110011001000;
   assign mem[14734] = 32'b11111000000111001101001011011000;
   assign mem[14735] = 32'b00000111010110111111110100011000;
   assign mem[14736] = 32'b11111011101100000011110011001000;
   assign mem[14737] = 32'b00001000011000001111100111110000;
   assign mem[14738] = 32'b00000010001011111100001111100000;
   assign mem[14739] = 32'b11110111010100001100101100100000;
   assign mem[14740] = 32'b11111100010000001110000010001100;
   assign mem[14741] = 32'b00000010101100110101100100110100;
   assign mem[14742] = 32'b00000111110000011110001011000000;
   assign mem[14743] = 32'b00000101001110000011011010001000;
   assign mem[14744] = 32'b11111010011010100001010100011000;
   assign mem[14745] = 32'b11111010010010110101011100111000;
   assign mem[14746] = 32'b00000001111101010101001001110010;
   assign mem[14747] = 32'b11110100010111000111100111110000;
   assign mem[14748] = 32'b00000001111100011110100101000110;
   assign mem[14749] = 32'b11110110000110111010111001100000;
   assign mem[14750] = 32'b00000001101010101110000000110000;
   assign mem[14751] = 32'b00000011001111100011101001111100;
   assign mem[14752] = 32'b11111110100101000001001101100010;
   assign mem[14753] = 32'b11111101001011010100101111001100;
   assign mem[14754] = 32'b11111110111101101011100110111100;
   assign mem[14755] = 32'b11111100101100100100111111110100;
   assign mem[14756] = 32'b00000001000101010110011110001010;
   assign mem[14757] = 32'b11110101010010111110111000000000;
   assign mem[14758] = 32'b11111110001101001110101111001110;
   assign mem[14759] = 32'b11110110100010101010110011010000;
   assign mem[14760] = 32'b00000010011010111110110101101000;
   assign mem[14761] = 32'b00000010001000100111001011111000;
   assign mem[14762] = 32'b00000100001011011000011100010000;
   assign mem[14763] = 32'b11111011101100101000011110111000;
   assign mem[14764] = 32'b11111011001001100010001000100000;
   assign mem[14765] = 32'b11111011111011011110100111000000;
   assign mem[14766] = 32'b00000100110101110010100001100000;
   assign mem[14767] = 32'b11111110100110011010111111001000;
   assign mem[14768] = 32'b00000000110100010011100101000000;
   assign mem[14769] = 32'b11111100001101000010110110110100;
   assign mem[14770] = 32'b00000100010101100001110010010000;
   assign mem[14771] = 32'b11110011000001011110100000100000;
   assign mem[14772] = 32'b11111111100111000011110111000100;
   assign mem[14773] = 32'b00000001111001101111011111110000;
   assign mem[14774] = 32'b11111101011001001010010101100000;
   assign mem[14775] = 32'b00000011111101111011110000000000;
   assign mem[14776] = 32'b11111110011000000100101011011000;
   assign mem[14777] = 32'b11111101011000110000101100100100;
   assign mem[14778] = 32'b00000010000001101011000011101000;
   assign mem[14779] = 32'b11111111010011010100010010101010;
   assign mem[14780] = 32'b00000000010101110111100011111100;
   assign mem[14781] = 32'b00000001011101111000001010111100;
   assign mem[14782] = 32'b11111000011001101111001101111000;
   assign mem[14783] = 32'b11111111011010111001101011110110;
   assign mem[14784] = 32'b11111111001010010111111010011000;
   assign mem[14785] = 32'b00000001011111111110000010010110;
   assign mem[14786] = 32'b00000001111011001000101000101110;
   assign mem[14787] = 32'b11111110111100011110110001000000;
   assign mem[14788] = 32'b00000000100011000101000101001000;
   assign mem[14789] = 32'b11111111000111110011001011010010;
   assign mem[14790] = 32'b00000100110010100101101110101000;
   assign mem[14791] = 32'b11110001001011011010111100000000;
   assign mem[14792] = 32'b00000001010000011000110001011100;
   assign mem[14793] = 32'b00000001111100011001111001011000;
   assign mem[14794] = 32'b11110110111010001100110111110000;
   assign mem[14795] = 32'b00000100100111100011001101000000;
   assign mem[14796] = 32'b00000010011011110000001111000100;
   assign mem[14797] = 32'b11111010101011010111011101111000;
   assign mem[14798] = 32'b00000011100001100110111011110100;
   assign mem[14799] = 32'b00000000001110000010000100001100;
   assign mem[14800] = 32'b00000101101101111001010001110000;
   assign mem[14801] = 32'b00000000010110010001001010001100;
   assign mem[14802] = 32'b00000100000111011000001001101000;
   assign mem[14803] = 32'b00000001101101011111001010010000;
   assign mem[14804] = 32'b11111010110111011001111001010000;
   assign mem[14805] = 32'b00000001011111011110000010000000;
   assign mem[14806] = 32'b00000010001101010000010101001000;
   assign mem[14807] = 32'b11101101101001000101000001100000;
   assign mem[14808] = 32'b11111100000101010111100111100000;
   assign mem[14809] = 32'b11111110111011101000011010010000;
   assign mem[14810] = 32'b11110111100011110110101111000000;
   assign mem[14811] = 32'b00000010010010001100101010101100;
   assign mem[14812] = 32'b11110000111010010000111001110000;
   assign mem[14813] = 32'b00000011110110111000010011010100;
   assign mem[14814] = 32'b11111110101110010010100101001100;
   assign mem[14815] = 32'b00000000100010010111010101010100;
   assign mem[14816] = 32'b11111010011010000110100100010000;
   assign mem[14817] = 32'b00000010011100001000111000011100;
   assign mem[14818] = 32'b11111101111000011110111110100000;
   assign mem[14819] = 32'b00000110001101111000100101101000;
   assign mem[14820] = 32'b00000000011101011101001001111011;
   assign mem[14821] = 32'b00000100111111111000111001100000;
   assign mem[14822] = 32'b11111101110011011010101001100100;
   assign mem[14823] = 32'b00000001010011100010011010101010;
   assign mem[14824] = 32'b11111110001101000110111110101010;
   assign mem[14825] = 32'b00000000110011100000111001110010;
   assign mem[14826] = 32'b11111110011000000011110111100000;
   assign mem[14827] = 32'b11110110010100111111111111010000;
   assign mem[14828] = 32'b11111111111010101010001001100101;
   assign mem[14829] = 32'b00000001100101101100110010100010;
   assign mem[14830] = 32'b00000000111111001001101000000100;
   assign mem[14831] = 32'b00000000010010011110111010101000;
   assign mem[14832] = 32'b00000101011100000100010001111000;
   assign mem[14833] = 32'b00000010001000011010110100000000;
   assign mem[14834] = 32'b00000010010000110011011010111000;
   assign mem[14835] = 32'b11111000111110001101001100001000;
   assign mem[14836] = 32'b00000001010101010010001110111010;
   assign mem[14837] = 32'b11111011010100110101010000111000;
   assign mem[14838] = 32'b11111110000010010111101000000000;
   assign mem[14839] = 32'b11111101011010000100101100101000;
   assign mem[14840] = 32'b11111111011000100110000110110000;
   assign mem[14841] = 32'b11111111010000110111001000101010;
   assign mem[14842] = 32'b00001110011011001110000001110000;
   assign mem[14843] = 32'b11111010010001110101001011010000;
   assign mem[14844] = 32'b11111110110011000101001011001010;
   assign mem[14845] = 32'b11111110011111001000110010000110;
   assign mem[14846] = 32'b00000011001100100100001111110100;
   assign mem[14847] = 32'b00000000100100110010110110101011;
   assign mem[14848] = 32'b11111011000101010111011011100000;
   assign mem[14849] = 32'b00000101000001110100001101001000;
   assign mem[14850] = 32'b11111101000111101111111111110100;
   assign mem[14851] = 32'b00000111110100110111010001010000;
   assign mem[14852] = 32'b00010011000011011110100010000000;
   assign mem[14853] = 32'b00000000011000001100011111010110;
   assign mem[14854] = 32'b11111110010100110000000110001100;
   assign mem[14855] = 32'b11111110010110001101100111111100;
   assign mem[14856] = 32'b11110110111100011011101010000000;
   assign mem[14857] = 32'b11111001110000100001000001111000;
   assign mem[14858] = 32'b11111101000000111010100000000100;
   assign mem[14859] = 32'b11111001101001100010010111010000;
   assign mem[14860] = 32'b00000000101001010101110111000001;
   assign mem[14861] = 32'b00000010101000000011000101110100;
   assign mem[14862] = 32'b00001010001000001001100011000000;
   assign mem[14863] = 32'b11110111011001110000101011100000;
   assign mem[14864] = 32'b11111010001001100010010101101000;
   assign mem[14865] = 32'b11111100100010111011011001101100;
   assign mem[14866] = 32'b00000100010110001010010011111000;
   assign mem[14867] = 32'b11111000010001000111010001001000;
   assign mem[14868] = 32'b00000100000101111101110101111000;
   assign mem[14869] = 32'b11111000100010101010001110011000;
   assign mem[14870] = 32'b11111001000010100010111011011000;
   assign mem[14871] = 32'b11110101011100011011100000100000;
   assign mem[14872] = 32'b11110001011010111100101100010000;
   assign mem[14873] = 32'b00000111011110110100110001011000;
   assign mem[14874] = 32'b00000000100100010110111010101101;
   assign mem[14875] = 32'b11111111110000010100010110001111;
   assign mem[14876] = 32'b11111000010001011010101100001000;
   assign mem[14877] = 32'b00000001111110111011001110000010;
   assign mem[14878] = 32'b00000000000111101011010100110010;
   assign mem[14879] = 32'b00000000101111111111100110101110;
   assign mem[14880] = 32'b00000010111001010100110000011000;
   assign mem[14881] = 32'b00000001101110100100110010110000;
   assign mem[14882] = 32'b00000000110010110001101110010000;
   assign mem[14883] = 32'b11111111001010110010011100011011;
   assign mem[14884] = 32'b11111001110101100000101110100000;
   assign mem[14885] = 32'b11111011000101111100100111000000;
   assign mem[14886] = 32'b00000001100111011100111110000100;
   assign mem[14887] = 32'b11111010010101111011001111111000;
   assign mem[14888] = 32'b11111101000110011011010011011100;
   assign mem[14889] = 32'b11111100110001100010001010110000;
   assign mem[14890] = 32'b11111000101111001110101101011000;
   assign mem[14891] = 32'b00000010101000011010000011000000;
   assign mem[14892] = 32'b00000100011011000111011000010000;
   assign mem[14893] = 32'b11111001001110011001101011110000;
   assign mem[14894] = 32'b00000010001000111111100001000100;
   assign mem[14895] = 32'b11111001111101111110010100110000;
   assign mem[14896] = 32'b11111100100010010111000000111100;
   assign mem[14897] = 32'b00000001111100001001001011110010;
   assign mem[14898] = 32'b11111010101000010000010101101000;
   assign mem[14899] = 32'b00000101001101000101110000100000;
   assign mem[14900] = 32'b00000100011001110001110001101000;
   assign mem[14901] = 32'b00000010011001000000111001000100;
   assign mem[14902] = 32'b00000101100111101101100100110000;
   assign mem[14903] = 32'b00000011010111010000011011111000;
   assign mem[14904] = 32'b11111100010001011000010001111100;
   assign mem[14905] = 32'b11111100010111001011110000101100;
   assign mem[14906] = 32'b00000001111110111100100010010010;
   assign mem[14907] = 32'b00000101111110000011110001011000;
   assign mem[14908] = 32'b00000001011111110111000000010110;
   assign mem[14909] = 32'b11110000001001011110100011010000;
   assign mem[14910] = 32'b00000101011111110000111111000000;
   assign mem[14911] = 32'b11101111100001001110000100000000;
   assign mem[14912] = 32'b00000001011011001110110000011100;
   assign mem[14913] = 32'b00000100011011011001101100011000;
   assign mem[14914] = 32'b11110001011010010100011101100000;
   assign mem[14915] = 32'b00000011000001011100111101100000;
   assign mem[14916] = 32'b00000011001100010111111111110100;
   assign mem[14917] = 32'b11111000110010000110010010111000;
   assign mem[14918] = 32'b00000100100111100000110111100000;
   assign mem[14919] = 32'b11111100111100011110111111011100;
   assign mem[14920] = 32'b11101010101101101010010001000000;
   assign mem[14921] = 32'b11111110110000110100111101010000;
   assign mem[14922] = 32'b11110111111000110111101111000000;
   assign mem[14923] = 32'b11111011111111001001001110011000;
   assign mem[14924] = 32'b00000111101010010101011000110000;
   assign mem[14925] = 32'b11111100100010100011011111001000;
   assign mem[14926] = 32'b11110010010100010010110111000000;
   assign mem[14927] = 32'b00001101100110011011100010110000;
   assign mem[14928] = 32'b11110111010001010100011100010000;
   assign mem[14929] = 32'b00001000111101101111000110110000;
   assign mem[14930] = 32'b00000011001011100010000100111100;
   assign mem[14931] = 32'b00000001001010110011100001100100;
   assign mem[14932] = 32'b00000011111001001000010110000000;
   assign mem[14933] = 32'b00000001010101000101010111011110;
   assign mem[14934] = 32'b11101110001010100000100001000000;
   assign mem[14935] = 32'b00000010111001110101101110000100;
   assign mem[14936] = 32'b11111111100110110100101001100011;
   assign mem[14937] = 32'b11110100011110111101001010110000;
   assign mem[14938] = 32'b00000011111000000010111011001000;
   assign mem[14939] = 32'b11111110111101110010100100010000;
   assign mem[14940] = 32'b00000001110100110010100011111100;
   assign mem[14941] = 32'b11101101110000011001110101000000;
   assign mem[14942] = 32'b11111111000010110001110111010000;
   assign mem[14943] = 32'b00000101001010010010000101001000;
   assign mem[14944] = 32'b11111001101001000111111101000000;
   assign mem[14945] = 32'b00000010111001111101111111001000;
   assign mem[14946] = 32'b00000001100011000010011000011110;
   assign mem[14947] = 32'b11111010101010100100011011100000;
   assign mem[14948] = 32'b00000101010100111101010011100000;
   assign mem[14949] = 32'b11111100100110110101100010110000;
   assign mem[14950] = 32'b11110001001000011111100011000000;
   assign mem[14951] = 32'b00000000111111100100011111111101;
   assign mem[14952] = 32'b00000010100111010001010101110100;
   assign mem[14953] = 32'b11111100000011100010010010101100;
   assign mem[14954] = 32'b00000001110010101011000110001100;
   assign mem[14955] = 32'b11111000110101110111100001101000;
   assign mem[14956] = 32'b11110111101101000001111000100000;
   assign mem[14957] = 32'b00000011111100011011111110011000;
   assign mem[14958] = 32'b11111110110110011001101111110010;
   assign mem[14959] = 32'b00000011010000110001001011110100;
   assign mem[14960] = 32'b11111011101101100111100010100000;
   assign mem[14961] = 32'b11111111010111100100111000011011;
   assign mem[14962] = 32'b00000101110001010010110101010000;
   assign mem[14963] = 32'b00000000010010100101110000110001;
   assign mem[14964] = 32'b00000010110000010000111100100000;
   assign mem[14965] = 32'b11111100000010100101101100011000;
   assign mem[14966] = 32'b11101111011100001110100100000000;
   assign mem[14967] = 32'b11111101001011100010101011011000;
   assign mem[14968] = 32'b11111110110000101001011101110000;
   assign mem[14969] = 32'b00000001010010111101101101010100;
   assign mem[14970] = 32'b11111100011011110000100111000000;
   assign mem[14971] = 32'b00000010100000101101010010010100;
   assign mem[14972] = 32'b11111000100010110100011101101000;
   assign mem[14973] = 32'b11111111010000110000011111010001;
   assign mem[14974] = 32'b00000000010000000001110100001101;
   assign mem[14975] = 32'b00000001011001001111111001111000;
   assign mem[14976] = 32'b11111110101000101011101111101000;
   assign mem[14977] = 32'b00000000100111111101110111000111;
   assign mem[14978] = 32'b11111111111101110010010011001101;
   assign mem[14979] = 32'b00000010111111011011011101010100;
   assign mem[14980] = 32'b11110110110111110000101101010000;
   assign mem[14981] = 32'b11111111100000001110011101001111;
   assign mem[14982] = 32'b11111000101101111101100010100000;
   assign mem[14983] = 32'b11111101001110011100000001100100;
   assign mem[14984] = 32'b00000011001101101110001110010100;
   assign mem[14985] = 32'b11111000110110101111000000101000;
   assign mem[14986] = 32'b11110101111011111000001110100000;
   assign mem[14987] = 32'b00000000110110011110111110011110;
   assign mem[14988] = 32'b00000010110101100000010001001100;
   assign mem[14989] = 32'b00000100111000111111001001110000;
   assign mem[14990] = 32'b00000111101111101101111111011000;
   assign mem[14991] = 32'b00000010000101001110111110000000;
   assign mem[14992] = 32'b11110110100101010110011000010000;
   assign mem[14993] = 32'b11111110110000000001000010100000;
   assign mem[14994] = 32'b11110101011000110000100001110000;
   assign mem[14995] = 32'b00000000001000000111011100111010;
   assign mem[14996] = 32'b00000111101010001110011000110000;
   assign mem[14997] = 32'b00000011011010101100011000000000;
   assign mem[14998] = 32'b11111010010001110111000001101000;
   assign mem[14999] = 32'b00000011010001110010100000001100;
   assign mem[15000] = 32'b00000101010010011000010100000000;
   assign mem[15001] = 32'b00000011100111010100110110111100;
   assign mem[15002] = 32'b00000011010010100101001011001000;
   assign mem[15003] = 32'b11111110011110110111110110111110;
   assign mem[15004] = 32'b11111000110000111111000100010000;
   assign mem[15005] = 32'b00000000010010010111110010111101;
   assign mem[15006] = 32'b00000100100100000011101100001000;
   assign mem[15007] = 32'b11111011110100001011011000101000;
   assign mem[15008] = 32'b00000011111101111001010001000100;
   assign mem[15009] = 32'b11111101001001010100101001010000;
   assign mem[15010] = 32'b00000101101001001100000111111000;
   assign mem[15011] = 32'b11110110110011010111011001000000;
   assign mem[15012] = 32'b00000101111010011011010101010000;
   assign mem[15013] = 32'b00000010001010000100101110010000;
   assign mem[15014] = 32'b11110110001100011111110001000000;
   assign mem[15015] = 32'b11111111010100111101101011000000;
   assign mem[15016] = 32'b00000100110000011011111010101000;
   assign mem[15017] = 32'b11110000101010010110000110100000;
   assign mem[15018] = 32'b00000001111110001110101011010100;
   assign mem[15019] = 32'b11110110101101000001011001110000;
   assign mem[15020] = 32'b11111010111100001110101101011000;
   assign mem[15021] = 32'b00000001001101110101001001101000;
   assign mem[15022] = 32'b11111001000111110101001100010000;
   assign mem[15023] = 32'b11111100100000111011101100100100;
   assign mem[15024] = 32'b00000101000100110100001100101000;
   assign mem[15025] = 32'b11111111001101011001011001001011;
   assign mem[15026] = 32'b11111100101100011101101100101100;
   assign mem[15027] = 32'b00000001001100110000010110110100;
   assign mem[15028] = 32'b00000000001110001111001011111001;
   assign mem[15029] = 32'b00000101001111000000111001001000;
   assign mem[15030] = 32'b00000100011101001100111011000000;
   assign mem[15031] = 32'b00000001110111000011000110110100;
   assign mem[15032] = 32'b00000011000001010010110010100100;
   assign mem[15033] = 32'b00000001011001111100010010100000;
   assign mem[15034] = 32'b11111100101111010000010011000100;
   assign mem[15035] = 32'b11111100100101000000111011100100;
   assign mem[15036] = 32'b11111110111101110011100101100010;
   assign mem[15037] = 32'b00000001110011000100000111010000;
   assign mem[15038] = 32'b11111110111010001110011111011100;
   assign mem[15039] = 32'b11111101110101111010001001010100;
   assign mem[15040] = 32'b00000111010000110101011011100000;
   assign mem[15041] = 32'b11110011000001001010110000110000;
   assign mem[15042] = 32'b00000010001111000001010000110100;
   assign mem[15043] = 32'b00000110001010100011101111100000;
   assign mem[15044] = 32'b11110100111011001010001001100000;
   assign mem[15045] = 32'b00000101100101011111011010000000;
   assign mem[15046] = 32'b11111100010110000011111001110100;
   assign mem[15047] = 32'b11111011110100000000001101101000;
   assign mem[15048] = 32'b11111010111011010101101101111000;
   assign mem[15049] = 32'b11111110111001001001111001100100;
   assign mem[15050] = 32'b11111101110101011111001100000000;
   assign mem[15051] = 32'b11110101011110110011010101000000;
   assign mem[15052] = 32'b11111100101011000101010010011000;
   assign mem[15053] = 32'b00001000000111110000110000000000;
   assign mem[15054] = 32'b00000000110001101101100111101001;
   assign mem[15055] = 32'b11111110100100010001000100110110;
   assign mem[15056] = 32'b00000100001111010100011001111000;
   assign mem[15057] = 32'b00000110010000001111101000010000;
   assign mem[15058] = 32'b11111101000100111000100110001000;
   assign mem[15059] = 32'b11111100100100101001000000100000;
   assign mem[15060] = 32'b00000001100000011100110010010000;
   assign mem[15061] = 32'b00000010110101100110001000011100;
   assign mem[15062] = 32'b00000100110100110001001000011000;
   assign mem[15063] = 32'b11111111000010011111000110010100;
   assign mem[15064] = 32'b11111110011011010010111101100100;
   assign mem[15065] = 32'b11111011001000100011111111110000;
   assign mem[15066] = 32'b00000010011001110110011011111100;
   assign mem[15067] = 32'b11111010000011010000010010111000;
   assign mem[15068] = 32'b00000001111110011100100010000000;
   assign mem[15069] = 32'b11110111010011110111101010000000;
   assign mem[15070] = 32'b00000100001011010110101100001000;
   assign mem[15071] = 32'b00000001111101001001100100100000;
   assign mem[15072] = 32'b11110110111001101000011001010000;
   assign mem[15073] = 32'b00000111000110111001011110111000;
   assign mem[15074] = 32'b11111111101101110110110010101011;
   assign mem[15075] = 32'b00000011100100011110100100010000;
   assign mem[15076] = 32'b00000001111000101010101110011110;
   assign mem[15077] = 32'b11111110111100010100011001001000;
   assign mem[15078] = 32'b00000100000101100000001000110000;
   assign mem[15079] = 32'b00000001000000101100011110101010;
   assign mem[15080] = 32'b00000100010101111101011011010000;
   assign mem[15081] = 32'b00000110000001001110011010010000;
   assign mem[15082] = 32'b00000110001100111100100001101000;
   assign mem[15083] = 32'b00000001100110110100000010101000;
   assign mem[15084] = 32'b11110010010110011100010100010000;
   assign mem[15085] = 32'b00000001011110111101011101000110;
   assign mem[15086] = 32'b00000010110001110011011001101000;
   assign mem[15087] = 32'b11111100010101110100100101110000;
   assign mem[15088] = 32'b00000011100010011000110101001000;
   assign mem[15089] = 32'b11101111101000001100011001000000;
   assign mem[15090] = 32'b11111000110000111001101101100000;
   assign mem[15091] = 32'b00001011001101000101011001010000;
   assign mem[15092] = 32'b00000110001100101101000100100000;
   assign mem[15093] = 32'b11111111011110000001111110011110;
   assign mem[15094] = 32'b00000101110110100101110111011000;
   assign mem[15095] = 32'b11111101001011001110001010110000;
   assign mem[15096] = 32'b11111111000001001000101001000001;
   assign mem[15097] = 32'b00000000001110011110100111011001;
   assign mem[15098] = 32'b00000001011011001101000111011010;
   assign mem[15099] = 32'b11110011010010111001101011000000;
   assign mem[15100] = 32'b00000001101101010011000010110010;
   assign mem[15101] = 32'b00001001001100011011100100110000;
   assign mem[15102] = 32'b00000011110101000100111101001000;
   assign mem[15103] = 32'b11110110010001000000000110100000;
   assign mem[15104] = 32'b00000000010100100100011011011111;
   assign mem[15105] = 32'b11111000111011010001000000011000;
   assign mem[15106] = 32'b00000101111110001100100010110000;
   assign mem[15107] = 32'b11111010101100111001011101001000;
   assign mem[15108] = 32'b00000010100111000110111101110100;
   assign mem[15109] = 32'b00000001101001110111100100011100;
   assign mem[15110] = 32'b00000011100101000111100010011100;
   assign mem[15111] = 32'b00000100010010000011101110000000;
   assign mem[15112] = 32'b00000010110100101001001111011100;
   assign mem[15113] = 32'b00000111010001000100101011010000;
   assign mem[15114] = 32'b11101101011000110110110011000000;
   assign mem[15115] = 32'b11111110100101111110101011011110;
   assign mem[15116] = 32'b00000101101000000000000001011000;
   assign mem[15117] = 32'b11110011111001101000111100100000;
   assign mem[15118] = 32'b00000000111110010010101111001111;
   assign mem[15119] = 32'b11111000001011011001010001100000;
   assign mem[15120] = 32'b11111100000111000111101001111100;
   assign mem[15121] = 32'b00000001101010101011001100110100;
   assign mem[15122] = 32'b00001001010111011101110010010000;
   assign mem[15123] = 32'b00000001000010000101101011100010;
   assign mem[15124] = 32'b11111111100111101111111000101000;
   assign mem[15125] = 32'b11110101110101110100010100100000;
   assign mem[15126] = 32'b00000011101011111100011100000100;
   assign mem[15127] = 32'b00000000011001010001001101001010;
   assign mem[15128] = 32'b11111001011011101000011110010000;
   assign mem[15129] = 32'b11111101110111011101000001001000;
   assign mem[15130] = 32'b00000011010110110001101111011000;
   assign mem[15131] = 32'b00000000010000000101100100010011;
   assign mem[15132] = 32'b00000001101001111000110100010110;
   assign mem[15133] = 32'b00000000010111010100000001001111;
   assign mem[15134] = 32'b11111101111000000011000101010000;
   assign mem[15135] = 32'b11111111100011001110010101100100;
   assign mem[15136] = 32'b00000100000100010000111111101000;
   assign mem[15137] = 32'b11111011000010110110111011100000;
   assign mem[15138] = 32'b11111010010100101110111111111000;
   assign mem[15139] = 32'b11111011111111011010010100001000;
   assign mem[15140] = 32'b00000010011101100010100101100000;
   assign mem[15141] = 32'b00000011001100010011110010011000;
   assign mem[15142] = 32'b00001000001001111011111011000000;
   assign mem[15143] = 32'b11111001110111101111100011100000;
   assign mem[15144] = 32'b11111100011111100001011101100100;
   assign mem[15145] = 32'b11111010000011010111011010101000;
   assign mem[15146] = 32'b00000111001001011111001111011000;
   assign mem[15147] = 32'b00000001100010110000011000111010;
   assign mem[15148] = 32'b11111100000010010111010001000100;
   assign mem[15149] = 32'b11110111100101101110111001010000;
   assign mem[15150] = 32'b11101101100000011101001001100000;
   assign mem[15151] = 32'b11111111111110000010010000110111;
   assign mem[15152] = 32'b11111111100011110110101011111110;
   assign mem[15153] = 32'b00000011110111100011001100011000;
   assign mem[15154] = 32'b11111010010011011010111010100000;
   assign mem[15155] = 32'b00001001000010010110100111000000;
   assign mem[15156] = 32'b11111100110110101010001000100000;
   assign mem[15157] = 32'b11111011101010101111110101000000;
   assign mem[15158] = 32'b00000110011001101010001000011000;
   assign mem[15159] = 32'b11111100010001000001100011111000;
   assign mem[15160] = 32'b11111111100100111110100011111010;
   assign mem[15161] = 32'b00000110110100011100101010100000;
   assign mem[15162] = 32'b00000110011001011011110110100000;
   assign mem[15163] = 32'b11101110101011011011111011000000;
   assign mem[15164] = 32'b11111111100101110001110011110111;
   assign mem[15165] = 32'b11110110000000111001001011000000;
   assign mem[15166] = 32'b00000011010101000000011111100000;
   assign mem[15167] = 32'b00000100010010100000110110100000;
   assign mem[15168] = 32'b11111110110000111111111011010010;
   assign mem[15169] = 32'b11111110000101101011100010111110;
   assign mem[15170] = 32'b11110100011011100111101011110000;
   assign mem[15171] = 32'b00000001011110111000110010001110;
   assign mem[15172] = 32'b00001001100110011100100110110000;
   assign mem[15173] = 32'b00001010010101010110101110010000;
   assign mem[15174] = 32'b11111000011000110100010100000000;
   assign mem[15175] = 32'b00001010011001101011000010110000;
   assign mem[15176] = 32'b11111010111000111010110010110000;
   assign mem[15177] = 32'b11110101011101111101011001110000;
   assign mem[15178] = 32'b00000011101000010111000011100000;
   assign mem[15179] = 32'b11101001110101101101111011000000;
   assign mem[15180] = 32'b11101101111000100110110100100000;
   assign mem[15181] = 32'b00010000011010110111110010000000;
   assign mem[15182] = 32'b00000000010000001000010000001010;
   assign mem[15183] = 32'b00000101110110100111000110011000;
   assign mem[15184] = 32'b00000110001100100001110101001000;
   assign mem[15185] = 32'b11110100001000000000111111000000;
   assign mem[15186] = 32'b11111001110010000000100010110000;
   assign mem[15187] = 32'b00000101101110010011011000000000;
   assign mem[15188] = 32'b11110011110001110000011011110000;
   assign mem[15189] = 32'b00000111011110010010110100101000;
   assign mem[15190] = 32'b00000010011101100000010011000000;
   assign mem[15191] = 32'b11111110011111011101110001011100;
   assign mem[15192] = 32'b11111100000011011111101001101100;
   assign mem[15193] = 32'b11111101001001110011110101100100;
   assign mem[15194] = 32'b11111110011100111000111000000100;
   assign mem[15195] = 32'b00000010011101000110000111100000;
   assign mem[15196] = 32'b11111110010101000001110010001100;
   assign mem[15197] = 32'b11111111100011000001101111010110;
   assign mem[15198] = 32'b00000000011110001100101101010111;
   assign mem[15199] = 32'b00000010000100000110000010101000;
   assign mem[15200] = 32'b00000001110010000001111010000100;
   assign mem[15201] = 32'b00000110011111100001000000111000;
   assign mem[15202] = 32'b00000101100010010111100001110000;
   assign mem[15203] = 32'b00000100110001000111001110110000;
   assign mem[15204] = 32'b11111101101100010000011011110100;
   assign mem[15205] = 32'b00000100100110100011010100001000;
   assign mem[15206] = 32'b00000011111100000100100000000100;
   assign mem[15207] = 32'b11111110000001110110001111010010;
   assign mem[15208] = 32'b11111100111001010011111111001100;
   assign mem[15209] = 32'b11111010010010010111001000000000;
   assign mem[15210] = 32'b00000101010000011000110110011000;
   assign mem[15211] = 32'b11111010000100010011100110011000;
   assign mem[15212] = 32'b11111110101100001111110000000010;
   assign mem[15213] = 32'b00000111111110100111111001110000;
   assign mem[15214] = 32'b11110100001110011100000110010000;
   assign mem[15215] = 32'b11111110010011111011010000110010;
   assign mem[15216] = 32'b00001000110000100001101010000000;
   assign mem[15217] = 32'b00000100100010001001110100000000;
   assign mem[15218] = 32'b00000001011000111010100110010010;
   assign mem[15219] = 32'b11111010010100011001111111010000;
   assign mem[15220] = 32'b11111101010100101111110000000100;
   assign mem[15221] = 32'b11111001101001001010001000110000;
   assign mem[15222] = 32'b11111111100001000101000110111101;
   assign mem[15223] = 32'b00000111100010000111000110111000;
   assign mem[15224] = 32'b11110011100000100100000010100000;
   assign mem[15225] = 32'b00000110111011011101000000101000;
   assign mem[15226] = 32'b00000011100100100000000110110000;
   assign mem[15227] = 32'b11110110111010101000101001110000;
   assign mem[15228] = 32'b00000110101100111011111111000000;
   assign mem[15229] = 32'b11111110100010000001010111101000;
   assign mem[15230] = 32'b11110001110010000011001001000000;
   assign mem[15231] = 32'b00000111111111110011011100101000;
   assign mem[15232] = 32'b00000101111111010000000011010000;
   assign mem[15233] = 32'b00000000110111111111101011001101;
   assign mem[15234] = 32'b00000101100010010001100010000000;
   assign mem[15235] = 32'b11110110111001000111001110110000;
   assign mem[15236] = 32'b11110110110010011111100000010000;
   assign mem[15237] = 32'b00001000001011011011001011010000;
   assign mem[15238] = 32'b11110101011110100110010111110000;
   assign mem[15239] = 32'b00001000100001010001110010100000;
   assign mem[15240] = 32'b00000010100011100100111010110000;
   assign mem[15241] = 32'b00000011101111110110111101010100;
   assign mem[15242] = 32'b00000011111110100010011111001000;
   assign mem[15243] = 32'b11111110110010110110111000001110;
   assign mem[15244] = 32'b00000001000000011100010101001010;
   assign mem[15245] = 32'b11111110001001111011010001100110;
   assign mem[15246] = 32'b00000011001011011111100100000100;
   assign mem[15247] = 32'b11110011111011101001101011100000;
   assign mem[15248] = 32'b00000000110110110001000111100011;
   assign mem[15249] = 32'b11111110000111011111010000100110;
   assign mem[15250] = 32'b00000101000000100110110000010000;
   assign mem[15251] = 32'b00000011000101011011110011000000;
   assign mem[15252] = 32'b00000100111011111010001110110000;
   assign mem[15253] = 32'b11111111000111010000010100011111;
   assign mem[15254] = 32'b11111010011001010001101010100000;
   assign mem[15255] = 32'b11111110101010101110100001100110;
   assign mem[15256] = 32'b00000110000000000011111000010000;
   assign mem[15257] = 32'b11110011000011111001100110010000;
   assign mem[15258] = 32'b00000001011111111010111011011000;
   assign mem[15259] = 32'b11111111110100101101110100011001;
   assign mem[15260] = 32'b00000011010011101001111000001100;
   assign mem[15261] = 32'b00000010010100111110110011011100;
   assign mem[15262] = 32'b00000000110010111000011100101010;
   assign mem[15263] = 32'b11111111110110001010000110000010;
   assign mem[15264] = 32'b11111001000101101110000011101000;
   assign mem[15265] = 32'b00000001101100011101110011110100;
   assign mem[15266] = 32'b00000000111111010110001100011101;
   assign mem[15267] = 32'b11110011111100000011110000100000;
   assign mem[15268] = 32'b00000001101100000011000011101100;
   assign mem[15269] = 32'b11111111110000111000110011001111;
   assign mem[15270] = 32'b00000010111101000001011011001100;
   assign mem[15271] = 32'b11110011111110110110101000100000;
   assign mem[15272] = 32'b11110101000001111111011011000000;
   assign mem[15273] = 32'b00000101010000000110010011111000;
   assign mem[15274] = 32'b11111011110010010111101011011000;
   assign mem[15275] = 32'b00001000110100011011001000000000;
   assign mem[15276] = 32'b00000001000101001101101101101000;
   assign mem[15277] = 32'b11111111001111000111110010101110;
   assign mem[15278] = 32'b00000101100110000011000110101000;
   assign mem[15279] = 32'b11111110111001010101001101101100;
   assign mem[15280] = 32'b11110101110100010010000111000000;
   assign mem[15281] = 32'b00000000001100101101011110011101;
   assign mem[15282] = 32'b11111001000000010100010100101000;
   assign mem[15283] = 32'b00000110010110111010110000000000;
   assign mem[15284] = 32'b11110111111011010000000111100000;
   assign mem[15285] = 32'b00001000101100000010100110010000;
   assign mem[15286] = 32'b00000100100101101100001010100000;
   assign mem[15287] = 32'b11111001110001010000001111101000;
   assign mem[15288] = 32'b00000110000101000111111000111000;
   assign mem[15289] = 32'b11110111001111000001001101000000;
   assign mem[15290] = 32'b11111110000111110010011010000010;
   assign mem[15291] = 32'b11111011111111111100110001000000;
   assign mem[15292] = 32'b00000011100110010000000010111100;
   assign mem[15293] = 32'b00000010100011110001111000011100;
   assign mem[15294] = 32'b11111101111001001100110100110100;
   assign mem[15295] = 32'b11111111111010101000011101001001;
   assign mem[15296] = 32'b00000001010111110011011111101000;
   assign mem[15297] = 32'b11111010100000000010101000100000;
   assign mem[15298] = 32'b11111000110111010110011000000000;
   assign mem[15299] = 32'b11111010001011010011011110011000;
   assign mem[15300] = 32'b11111111101100011001010110100110;
   assign mem[15301] = 32'b11111010000111100111100011010000;
   assign mem[15302] = 32'b00000000010010010101010010100011;
   assign mem[15303] = 32'b00001000110000110000110011100000;
   assign mem[15304] = 32'b11110001000000011010010010110000;
   assign mem[15305] = 32'b00000110011111110100100001101000;
   assign mem[15306] = 32'b11111110000011101001001001101100;
   assign mem[15307] = 32'b11110000000001101111011110010000;
   assign mem[15308] = 32'b00000010010111000010110100100100;
   assign mem[15309] = 32'b11111000010000001100011011101000;
   assign mem[15310] = 32'b11110110111011101111101100110000;
   assign mem[15311] = 32'b00000000110100011011111001011110;
   assign mem[15312] = 32'b00000011100101011111100011100100;
   assign mem[15313] = 32'b00000011110100000101010100110000;
   assign mem[15314] = 32'b11110111011100001010001010000000;
   assign mem[15315] = 32'b00000110011100100101110001000000;
   assign mem[15316] = 32'b00000011100010001111001100010000;
   assign mem[15317] = 32'b11110000101010110000010110000000;
   assign mem[15318] = 32'b00001000101010000010101001100000;
   assign mem[15319] = 32'b11110111011011110010101010110000;
   assign mem[15320] = 32'b00000100101001011100100101110000;
   assign mem[15321] = 32'b00000011110100101110101001111100;
   assign mem[15322] = 32'b00000111011010010111010011101000;
   assign mem[15323] = 32'b00001001111010011011010101000000;
   assign mem[15324] = 32'b11101100000100011001010100000000;
   assign mem[15325] = 32'b00000101100100101101101001101000;
   assign mem[15326] = 32'b00000010110101110011110101101100;
   assign mem[15327] = 32'b11111011110001101100101111111000;
   assign mem[15328] = 32'b00000010110001000110100111101100;
   assign mem[15329] = 32'b11110001111001110100001010110000;
   assign mem[15330] = 32'b00000110001001110101100010000000;
   assign mem[15331] = 32'b11110011010001100101000101110000;
   assign mem[15332] = 32'b11111100000000011100010100111000;
   assign mem[15333] = 32'b00000101000011101011001110000000;
   assign mem[15334] = 32'b11110110100101101001111100110000;
   assign mem[15335] = 32'b00000010101110111010111101010000;
   assign mem[15336] = 32'b11111111110001000010010100101100;
   assign mem[15337] = 32'b00001110011111101010011110000000;
   assign mem[15338] = 32'b11111011101100001111001100101000;
   assign mem[15339] = 32'b11111011011101100111101100100000;
   assign mem[15340] = 32'b11110000011111010000000110110000;
   assign mem[15341] = 32'b00000100101000011001000000111000;
   assign mem[15342] = 32'b11110111101111100111111100110000;
   assign mem[15343] = 32'b11111001101101110001001011010000;
   assign mem[15344] = 32'b00000100000001011101110110110000;
   assign mem[15345] = 32'b11110101001011010011111111110000;
   assign mem[15346] = 32'b11101101111110011010100001000000;
   assign mem[15347] = 32'b00001001000011000100010010010000;
   assign mem[15348] = 32'b11101101010000011101110000000000;
   assign mem[15349] = 32'b00001000000100011011111101010000;
   assign mem[15350] = 32'b00000000110001110100111100111100;
   assign mem[15351] = 32'b11110110110001101011110101110000;
   assign mem[15352] = 32'b11110110110000101110101110110000;
   assign mem[15353] = 32'b00001000000010001001100011110000;
   assign mem[15354] = 32'b11111110011011011110110001001000;
   assign mem[15355] = 32'b11111110100011101100010001011010;
   assign mem[15356] = 32'b11111101101101000110100101000000;
   assign mem[15357] = 32'b11111110110100110110111111001010;
   assign mem[15358] = 32'b11111110011111000001011011100010;
   assign mem[15359] = 32'b11111110111101010100011100010000;
   assign mem[15360] = 32'b00001000001001010101101011110000;
   assign mem[15361] = 32'b11111011011001101101110001011000;
   assign mem[15362] = 32'b00000101001000110001010000110000;
   assign mem[15363] = 32'b11111010010111000010010101001000;
   assign mem[15364] = 32'b11101111111011111111101101100000;
   assign mem[15365] = 32'b00000101110100111101110011000000;
   assign mem[15366] = 32'b11111110100111010010000111101100;
   assign mem[15367] = 32'b00000010111111111101111101100100;
   assign mem[15368] = 32'b00000001011111100110010000100000;
   assign mem[15369] = 32'b11111111101111110010011000111010;
   assign mem[15370] = 32'b11101001100001011011011001000000;
   assign mem[15371] = 32'b00000110111110110100011111110000;
   assign mem[15372] = 32'b00000100010111100111001100101000;
   assign mem[15373] = 32'b00000010000010000101001000000000;
   assign mem[15374] = 32'b11111011110100110110101001000000;
   assign mem[15375] = 32'b11111110011110110011010010010000;
   assign mem[15376] = 32'b11111010101100110101001000000000;
   assign mem[15377] = 32'b11111010001100110011111000111000;
   assign mem[15378] = 32'b00000011111101100001011000111000;
   assign mem[15379] = 32'b00000000110001001011111011000100;
   assign mem[15380] = 32'b11101111001101111110110001100000;
   assign mem[15381] = 32'b00001001000010111011011001110000;
   assign mem[15382] = 32'b00001100000010010101111110010000;
   assign mem[15383] = 32'b11111011110111001001000110100000;
   assign mem[15384] = 32'b00000100110011010100011000001000;
   assign mem[15385] = 32'b11110101001010111001000001110000;
   assign mem[15386] = 32'b11111101001000101011001000110000;
   assign mem[15387] = 32'b11110011001101111000100110110000;
   assign mem[15388] = 32'b11111110000110101011101000001100;
   assign mem[15389] = 32'b00000000001000000100010110001110;
   assign mem[15390] = 32'b00000001101000001101010100001110;
   assign mem[15391] = 32'b00000110101011011111100100111000;
   assign mem[15392] = 32'b00000111000100000001011010000000;
   assign mem[15393] = 32'b11110110010110011000010010110000;
   assign mem[15394] = 32'b00000101000111001101000100010000;
   assign mem[15395] = 32'b11111000001110000011000101010000;
   assign mem[15396] = 32'b00000100011101111011011000100000;
   assign mem[15397] = 32'b00000001111010010000011101001010;
   assign mem[15398] = 32'b11110011000110111110101001110000;
   assign mem[15399] = 32'b11110110010010000000000111010000;
   assign mem[15400] = 32'b00000011111100110111011110010100;
   assign mem[15401] = 32'b11111111101000001001101110011000;
   assign mem[15402] = 32'b00000001110100011111111110100000;
   assign mem[15403] = 32'b11111011100101000111000011110000;
   assign mem[15404] = 32'b00000010101110001001111011110100;
   assign mem[15405] = 32'b11111011011010011001101111011000;
   assign mem[15406] = 32'b00000011101100111001111111000100;
   assign mem[15407] = 32'b11111111000100101000010011100111;
   assign mem[15408] = 32'b11111101110001110111101101010000;
   assign mem[15409] = 32'b11110111010010001010110100010000;
   assign mem[15410] = 32'b00000011110111000100100111010000;
   assign mem[15411] = 32'b11110110111000000101001001100000;
   assign mem[15412] = 32'b11110110111101111010001011100000;
   assign mem[15413] = 32'b00000110000101110101001010000000;
   assign mem[15414] = 32'b11111100100100010010110010011000;
   assign mem[15415] = 32'b00000110000010111010001000011000;
   assign mem[15416] = 32'b11110111111010100001100001000000;
   assign mem[15417] = 32'b11111101110101000110100101101000;
   assign mem[15418] = 32'b00000110000010010001010011001000;
   assign mem[15419] = 32'b11111011110001010010101010100000;
   assign mem[15420] = 32'b00000000100010001011010011100101;
   assign mem[15421] = 32'b11111101110111001100011001010100;
   assign mem[15422] = 32'b11111110001111000000011001101010;
   assign mem[15423] = 32'b00000001000110011011101101011010;
   assign mem[15424] = 32'b11111110101101110000101100111000;
   assign mem[15425] = 32'b11111111101000111001010111010100;
   assign mem[15426] = 32'b00000000100010110000101010111000;
   assign mem[15427] = 32'b11111111100100011010101101000011;
   assign mem[15428] = 32'b11111110101101011010000010011010;
   assign mem[15429] = 32'b11111011011111010101100001011000;
   assign mem[15430] = 32'b00000111001011000000110101001000;
   assign mem[15431] = 32'b11111001011111100001000011100000;
   assign mem[15432] = 32'b11111001101101011111001011011000;
   assign mem[15433] = 32'b00000010000000110100001011000100;
   assign mem[15434] = 32'b11110011100001010100100101100000;
   assign mem[15435] = 32'b00000000011100000010111011000001;
   assign mem[15436] = 32'b00000000001101010010110000011101;
   assign mem[15437] = 32'b11111110001000110101010000111110;
   assign mem[15438] = 32'b11111111111100101000100011010100;
   assign mem[15439] = 32'b11111100001011100100100100000000;
   assign mem[15440] = 32'b11111111110100000000000000111111;
   assign mem[15441] = 32'b00000111000001111100110001101000;
   assign mem[15442] = 32'b00010011001100111111011100000000;
   assign mem[15443] = 32'b11110001111001001110001010000000;
   assign mem[15444] = 32'b00001000110000011101100001010000;
   assign mem[15445] = 32'b11111000101001100100110000101000;
   assign mem[15446] = 32'b11101100110110100110001111100000;
   assign mem[15447] = 32'b11110011000100011101111000000000;
   assign mem[15448] = 32'b11110100101110100101010011010000;
   assign mem[15449] = 32'b00000110011111001010001111000000;
   assign mem[15450] = 32'b00001000001110001010100100100000;
   assign mem[15451] = 32'b11110001001110111100110011100000;
   assign mem[15452] = 32'b11111000000011010010111000100000;
   assign mem[15453] = 32'b00001000000000100010110111100000;
   assign mem[15454] = 32'b11111011100001100010100101110000;
   assign mem[15455] = 32'b11111111111110011100111101111000;
   assign mem[15456] = 32'b00000110000110111101111111000000;
   assign mem[15457] = 32'b11111100010011100101110001100000;
   assign mem[15458] = 32'b00000000000110111010101000001011;
   assign mem[15459] = 32'b11111011101100101001011000000000;
   assign mem[15460] = 32'b00000001100011101111100100000100;
   assign mem[15461] = 32'b00000011101100101010100000010100;
   assign mem[15462] = 32'b00001010111100010111101000000000;
   assign mem[15463] = 32'b11111000000010110111111000100000;
   assign mem[15464] = 32'b00000010011011011000110010011100;
   assign mem[15465] = 32'b11111011010111101000000111000000;
   assign mem[15466] = 32'b11111011011110000001110110000000;
   assign mem[15467] = 32'b11110101100001010110101111100000;
   assign mem[15468] = 32'b11111110011101100101110110111100;
   assign mem[15469] = 32'b00000001011110110111110111001110;
   assign mem[15470] = 32'b11110110000000101011111001010000;
   assign mem[15471] = 32'b00000110110010111010101101001000;
   assign mem[15472] = 32'b00001101011101010011110001010000;
   assign mem[15473] = 32'b11110000110111100010001001100000;
   assign mem[15474] = 32'b00001000100001101110000001010000;
   assign mem[15475] = 32'b11111011110011100000011011010000;
   assign mem[15476] = 32'b11111100100001000010011111011000;
   assign mem[15477] = 32'b11111010111010000011000001101000;
   assign mem[15478] = 32'b11110111101101100101101100010000;
   assign mem[15479] = 32'b00000110001011010010110111101000;
   assign mem[15480] = 32'b11110011000001011010100001010000;
   assign mem[15481] = 32'b11111000000111110010000010110000;
   assign mem[15482] = 32'b00011011000010001001100101100000;
   assign mem[15483] = 32'b11110111010101100111111010010000;
   assign mem[15484] = 32'b00000100101011010001101001010000;
   assign mem[15485] = 32'b11110100000011110110110000100000;
   assign mem[15486] = 32'b00000000101100001001010011111110;
   assign mem[15487] = 32'b11110101101111100001111100010000;
   assign mem[15488] = 32'b11110010110000010111100001000000;
   assign mem[15489] = 32'b00000110111110011001101011111000;
   assign mem[15490] = 32'b11101000101101000010111010000000;
   assign mem[15491] = 32'b00000010111001101011110100110000;
   assign mem[15492] = 32'b00010100100101100100100011100000;
   assign mem[15493] = 32'b11111000001101110011101010100000;
   assign mem[15494] = 32'b00001010110100001011111101010000;
   assign mem[15495] = 32'b11110100101111111100000011000000;
   assign mem[15496] = 32'b11110100010000100110001011110000;
   assign mem[15497] = 32'b11110100110000000010111010110000;
   assign mem[15498] = 32'b11110110110111001011100000110000;
   assign mem[15499] = 32'b11111111110001101000111010001011;
   assign mem[15500] = 32'b11111000011110000011000101101000;
   assign mem[15501] = 32'b00000101111101000101111010101000;
   assign mem[15502] = 32'b00001111011111011000010010010000;
   assign mem[15503] = 32'b11111100101011111100101010101000;
   assign mem[15504] = 32'b00000100001110011100010100100000;
   assign mem[15505] = 32'b11111001111000111001111000110000;
   assign mem[15506] = 32'b11111101100111011111011111010000;
   assign mem[15507] = 32'b11111011001001001001111100110000;
   assign mem[15508] = 32'b11110101111111101100101011110000;
   assign mem[15509] = 32'b00000001000001000011010010011100;
   assign mem[15510] = 32'b11111111110100011011111000010001;
   assign mem[15511] = 32'b11111010000001001001110010011000;
   assign mem[15512] = 32'b11110000000011101101001110100000;
   assign mem[15513] = 32'b00000110100000001101100000100000;
   assign mem[15514] = 32'b11111100001110101100001100001100;
   assign mem[15515] = 32'b11111111111111101100000000000111;
   assign mem[15516] = 32'b11111011111001101000111110100000;
   assign mem[15517] = 32'b11111001001100111000101111111000;
   assign mem[15518] = 32'b00001000100010000001110010100000;
   assign mem[15519] = 32'b11111001110111011010110010111000;
   assign mem[15520] = 32'b00000001100011010011100111110100;
   assign mem[15521] = 32'b00000011110011111101110011110000;
   assign mem[15522] = 32'b00001000110111111110111010100000;
   assign mem[15523] = 32'b11111010000111111111010001111000;
   assign mem[15524] = 32'b00000110010111111001010000011000;
   assign mem[15525] = 32'b11111100111000001101010101011000;
   assign mem[15526] = 32'b00000011110110000100010111000100;
   assign mem[15527] = 32'b11110010101011111011100010110000;
   assign mem[15528] = 32'b00000000001000001110000111000001;
   assign mem[15529] = 32'b11110110011000101101101101010000;
   assign mem[15530] = 32'b11111111010110001001000011000001;
   assign mem[15531] = 32'b11111110101110101100111001001010;
   assign mem[15532] = 32'b00000011000011111100010111100100;
   assign mem[15533] = 32'b11110110110100010111011101110000;
   assign mem[15534] = 32'b00001101011110110100000101110000;
   assign mem[15535] = 32'b11111000111111000010111111100000;
   assign mem[15536] = 32'b11111110101101100101011000100100;
   assign mem[15537] = 32'b11110000001110111111111110100000;
   assign mem[15538] = 32'b00000011001010110101110101101000;
   assign mem[15539] = 32'b00000110011000001011000110110000;
   assign mem[15540] = 32'b00001000111000101000001011100000;
   assign mem[15541] = 32'b00000000010101111011100010010010;
   assign mem[15542] = 32'b00000111010011111100000111101000;
   assign mem[15543] = 32'b11111011100101110101011010011000;
   assign mem[15544] = 32'b00000001101100101111010010101100;
   assign mem[15545] = 32'b11110010100100011101001110010000;
   assign mem[15546] = 32'b00000001010111001010101101001100;
   assign mem[15547] = 32'b00000010101001111000101111011000;
   assign mem[15548] = 32'b11111111111110001001000001000110;
   assign mem[15549] = 32'b11111000101010111000011110110000;
   assign mem[15550] = 32'b00001111011011000101010101000000;
   assign mem[15551] = 32'b11111111101000111100000011001100;
   assign mem[15552] = 32'b11111101111101000111101011110000;
   assign mem[15553] = 32'b00000101111010010010000110001000;
   assign mem[15554] = 32'b11111101101101000001001010000100;
   assign mem[15555] = 32'b11111111010011110011000111000000;
   assign mem[15556] = 32'b00000100000000001001111110100000;
   assign mem[15557] = 32'b11110111100011010011010110000000;
   assign mem[15558] = 32'b00000010010011111011010000101100;
   assign mem[15559] = 32'b11101100110011001100101000100000;
   assign mem[15560] = 32'b11101110111100110011000111100000;
   assign mem[15561] = 32'b11111110110011110111000110101010;
   assign mem[15562] = 32'b00000000110000100001101100000000;
   assign mem[15563] = 32'b11111101100111101000000100011000;
   assign mem[15564] = 32'b00001101100110110100010101110000;
   assign mem[15565] = 32'b00000000011000001000001000001100;
   assign mem[15566] = 32'b11101101001001110000110100000000;
   assign mem[15567] = 32'b11111010001110100010111000100000;
   assign mem[15568] = 32'b00000010100010110010101111101100;
   assign mem[15569] = 32'b00001001000111101110101101100000;
   assign mem[15570] = 32'b11111110000100101110110100111100;
   assign mem[15571] = 32'b00000000010111111110001111111110;
   assign mem[15572] = 32'b00001101000000100010010111010000;
   assign mem[15573] = 32'b00000000000111100000011110010110;
   assign mem[15574] = 32'b00000110000101111000100010100000;
   assign mem[15575] = 32'b00000001111101100000001101101110;
   assign mem[15576] = 32'b00000001000000001100100000110110;
   assign mem[15577] = 32'b11110011001000110101010000000000;
   assign mem[15578] = 32'b00000000101010000101010000000000;
   assign mem[15579] = 32'b11110100110010110000000000010000;
   assign mem[15580] = 32'b00000100110000011000001111111000;
   assign mem[15581] = 32'b11111000011100100010010100011000;
   assign mem[15582] = 32'b11110101010110011000010010010000;
   assign mem[15583] = 32'b00000101111000100011110011101000;
   assign mem[15584] = 32'b11110010101001110000010110000000;
   assign mem[15585] = 32'b00000011010001000100101000101000;
   assign mem[15586] = 32'b00000010011000111010110010111000;
   assign mem[15587] = 32'b11111100011010100010110101100000;
   assign mem[15588] = 32'b00000011110100101010110001111100;
   assign mem[15589] = 32'b11111011101101100100000111011000;
   assign mem[15590] = 32'b11110010111100110111010110000000;
   assign mem[15591] = 32'b00001000110111010110000100000000;
   assign mem[15592] = 32'b00000000011011110101110100010011;
   assign mem[15593] = 32'b11111101001001111100111011111000;
   assign mem[15594] = 32'b00000010101011001011011101010100;
   assign mem[15595] = 32'b11111011110001111001011100010000;
   assign mem[15596] = 32'b11110011001010001110011000000000;
   assign mem[15597] = 32'b11111100000111110000100110110100;
   assign mem[15598] = 32'b11111111111101010101011010110001;
   assign mem[15599] = 32'b00001001011101011100000001000000;
   assign mem[15600] = 32'b11101110110001111011110100000000;
   assign mem[15601] = 32'b11111100110111011100110001111000;
   assign mem[15602] = 32'b00000010001110101001010100011100;
   assign mem[15603] = 32'b00000000111101011000101100000001;
   assign mem[15604] = 32'b00000001100100111110000010111010;
   assign mem[15605] = 32'b11111011011111111010001101001000;
   assign mem[15606] = 32'b11111010011001011011110100111000;
   assign mem[15607] = 32'b11111000000000111110101001001000;
   assign mem[15608] = 32'b00000001010011010010011100101010;
   assign mem[15609] = 32'b00001001100101100010100010000000;
   assign mem[15610] = 32'b11111110011000011000111111111010;
   assign mem[15611] = 32'b11111110011101100101100000000010;
   assign mem[15612] = 32'b11111101010011101000111100110100;
   assign mem[15613] = 32'b00000100000010000101100110001000;
   assign mem[15614] = 32'b00000010100111010101011011001000;
   assign mem[15615] = 32'b11111111001100101000100000011000;
   assign mem[15616] = 32'b11111111101011110110000011110110;
   assign mem[15617] = 32'b00000000001011100011011101101000;
   assign mem[15618] = 32'b11111111001100100100101110000000;
   assign mem[15619] = 32'b11111101001110111110000000001100;
   assign mem[15620] = 32'b11111010100010011001001100001000;
   assign mem[15621] = 32'b11111011111101111111010111011000;
   assign mem[15622] = 32'b00000001011110110001110010011110;
   assign mem[15623] = 32'b11111110111111101100001011001100;
   assign mem[15624] = 32'b00000010101000000010011000111000;
   assign mem[15625] = 32'b11111010011100110010100000011000;
   assign mem[15626] = 32'b11111010011000001000111111010000;
   assign mem[15627] = 32'b00000101111001000001011100000000;
   assign mem[15628] = 32'b11111101111111010101100000010100;
   assign mem[15629] = 32'b00000011100101000101001111100000;
   assign mem[15630] = 32'b00001011101110110000101001000000;
   assign mem[15631] = 32'b11101100000111111000100111100000;
   assign mem[15632] = 32'b11110101100111101100011110100000;
   assign mem[15633] = 32'b00000110111101011110111100010000;
   assign mem[15634] = 32'b00000001000111101011000011000000;
   assign mem[15635] = 32'b00000010001111011111010110100100;
   assign mem[15636] = 32'b00001000101001110011110101110000;
   assign mem[15637] = 32'b00000111011101010001011001101000;
   assign mem[15638] = 32'b11111110100110101110010101001100;
   assign mem[15639] = 32'b11111100011111011101001011100100;
   assign mem[15640] = 32'b11111000011000011010111100000000;
   assign mem[15641] = 32'b00000000000000001110010000111011;
   assign mem[15642] = 32'b00001001110000110010010010010000;
   assign mem[15643] = 32'b11111011101100100010100100001000;
   assign mem[15644] = 32'b00000000111111001001000011011001;
   assign mem[15645] = 32'b11111110000110101110100000111010;
   assign mem[15646] = 32'b00000101010001110100011010101000;
   assign mem[15647] = 32'b11111000101100011011011110101000;
   assign mem[15648] = 32'b00000101101101010001111000101000;
   assign mem[15649] = 32'b11111101010011010111000101011000;
   assign mem[15650] = 32'b00000010010110001001001111100100;
   assign mem[15651] = 32'b00000111101101100110110101011000;
   assign mem[15652] = 32'b00010101101000110110101100100000;
   assign mem[15653] = 32'b11101110101111101101010010100000;
   assign mem[15654] = 32'b00000010010101111011001111101100;
   assign mem[15655] = 32'b11111111000001011110000111000010;
   assign mem[15656] = 32'b11110011111010000000110100100000;
   assign mem[15657] = 32'b11101111100011101000100011000000;
   assign mem[15658] = 32'b11111000011011111011010111101000;
   assign mem[15659] = 32'b11111000001001001110000001010000;
   assign mem[15660] = 32'b11110101011100000100101111100000;
   assign mem[15661] = 32'b11111011110111010000000000101000;
   assign mem[15662] = 32'b11101110100100111111000110100000;
   assign mem[15663] = 32'b00000011110111111010110111010100;
   assign mem[15664] = 32'b11111111111011111001010110010111;
   assign mem[15665] = 32'b11111111011011110110010001001110;
   assign mem[15666] = 32'b11111111110100111101001001010100;
   assign mem[15667] = 32'b00000011101011010010001000101100;
   assign mem[15668] = 32'b00000011000000101100110001100000;
   assign mem[15669] = 32'b00000000010111100011100000111100;
   assign mem[15670] = 32'b00000000100101010011110011100010;
   assign mem[15671] = 32'b00000101101000101111011110010000;
   assign mem[15672] = 32'b00000110111100110111010101010000;
   assign mem[15673] = 32'b11111010000001101101100011110000;
   assign mem[15674] = 32'b00000111101001000101001010000000;
   assign mem[15675] = 32'b11110110010011100010000101010000;
   assign mem[15676] = 32'b11111101000000000101001001100000;
   assign mem[15677] = 32'b00000001111000010000111010000000;
   assign mem[15678] = 32'b00000001001101101000010110001000;
   assign mem[15679] = 32'b11110100010011011001011000110000;
   assign mem[15680] = 32'b00000111011001100000011100010000;
   assign mem[15681] = 32'b11110001011111101111011100110000;
   assign mem[15682] = 32'b11110101111110010111011111100000;
   assign mem[15683] = 32'b00000110101101011001001000110000;
   assign mem[15684] = 32'b11101110111101000111110110000000;
   assign mem[15685] = 32'b00000111110000101101101000011000;
   assign mem[15686] = 32'b00000011101110010011001011010000;
   assign mem[15687] = 32'b11111011000101110100111011001000;
   assign mem[15688] = 32'b00000100100111101010100011011000;
   assign mem[15689] = 32'b11110111010111011010111111110000;
   assign mem[15690] = 32'b00000000010110110100011111100100;
   assign mem[15691] = 32'b11111100101011000100101100001100;
   assign mem[15692] = 32'b11110011101011000010011010110000;
   assign mem[15693] = 32'b00000100110000001111000111011000;
   assign mem[15694] = 32'b11111011110111001100100101010000;
   assign mem[15695] = 32'b00000100000010101001000110001000;
   assign mem[15696] = 32'b11111100011110101011101111000100;
   assign mem[15697] = 32'b11111100010101101101110000110100;
   assign mem[15698] = 32'b11111111010111010110010100010100;
   assign mem[15699] = 32'b00000011101111110100000100101100;
   assign mem[15700] = 32'b11111111010111001011001100101000;
   assign mem[15701] = 32'b00000111110111001011010011101000;
   assign mem[15702] = 32'b00000110011000101100000011111000;
   assign mem[15703] = 32'b11111010001101110101101111011000;
   assign mem[15704] = 32'b11111111100111111011100010000001;
   assign mem[15705] = 32'b11110110111000101010001010100000;
   assign mem[15706] = 32'b00000000000001000101100110101101;
   assign mem[15707] = 32'b11111100011111100110010000101000;
   assign mem[15708] = 32'b11111100011011100110101001110000;
   assign mem[15709] = 32'b11111101010010000100100111110000;
   assign mem[15710] = 32'b00000011011001101001100000001000;
   assign mem[15711] = 32'b11111011100011011001111101011000;
   assign mem[15712] = 32'b11111010011011110001000010110000;
   assign mem[15713] = 32'b00000001000100111110100100000000;
   assign mem[15714] = 32'b11111101100011001010001010001100;
   assign mem[15715] = 32'b00000010101101001111011000011100;
   assign mem[15716] = 32'b00000010010101001001000010010000;
   assign mem[15717] = 32'b11111111001000011001110101001010;
   assign mem[15718] = 32'b00000000110001011101101110111100;
   assign mem[15719] = 32'b11111100111101011111100111010100;
   assign mem[15720] = 32'b00000010100111011001101000010100;
   assign mem[15721] = 32'b00001100000111011101110010100000;
   assign mem[15722] = 32'b00010100000110000010011101000000;
   assign mem[15723] = 32'b11110110000110110110001100000000;
   assign mem[15724] = 32'b00000000111001100110101100110110;
   assign mem[15725] = 32'b11110000111101110011001000100000;
   assign mem[15726] = 32'b11111010110000101010110000001000;
   assign mem[15727] = 32'b11111011111011110000001010101000;
   assign mem[15728] = 32'b11111001100111000111011100110000;
   assign mem[15729] = 32'b11111100010011111000011001001100;
   assign mem[15730] = 32'b11110001000110100011010111000000;
   assign mem[15731] = 32'b00001001000101100110010001100000;
   assign mem[15732] = 32'b00001010000101110101001000100000;
   assign mem[15733] = 32'b11110110101100101101100100010000;
   assign mem[15734] = 32'b00000101010111110110110010011000;
   assign mem[15735] = 32'b11110110111100110011111110110000;
   assign mem[15736] = 32'b11111001001001000010111010010000;
   assign mem[15737] = 32'b11110101111010100001111010010000;
   assign mem[15738] = 32'b11111100001111111000000001011100;
   assign mem[15739] = 32'b00000000110100011001011000110010;
   assign mem[15740] = 32'b11110011100001101010110101100000;
   assign mem[15741] = 32'b00001101011111111101111011100000;
   assign mem[15742] = 32'b00001110010011000111100100010000;
   assign mem[15743] = 32'b11111010111110001001100100001000;
   assign mem[15744] = 32'b00001000110010000111011110000000;
   assign mem[15745] = 32'b11111001000010110010001001011000;
   assign mem[15746] = 32'b11111001000111100000101010000000;
   assign mem[15747] = 32'b11111101110110101110111110001000;
   assign mem[15748] = 32'b11110111110100101010001111110000;
   assign mem[15749] = 32'b00000011111010001011110011101000;
   assign mem[15750] = 32'b00000110101111100100110101110000;
   assign mem[15751] = 32'b00001000001000110001110000100000;
   assign mem[15752] = 32'b00000101001111110110111000010000;
   assign mem[15753] = 32'b11111000011000000000001111100000;
   assign mem[15754] = 32'b00000000010010000011110001100010;
   assign mem[15755] = 32'b11111000100011101110000011111000;
   assign mem[15756] = 32'b00001001010001000000111001110000;
   assign mem[15757] = 32'b11111010101111100000011100110000;
   assign mem[15758] = 32'b11111111000100100110100110101010;
   assign mem[15759] = 32'b11110111111110110101000010000000;
   assign mem[15760] = 32'b11111111111001100100011100100000;
   assign mem[15761] = 32'b00000010000010000001011100100100;
   assign mem[15762] = 32'b00000111011001000101000001101000;
   assign mem[15763] = 32'b11111100110111010011111101011100;
   assign mem[15764] = 32'b00000011100011101001101110001000;
   assign mem[15765] = 32'b11110110001011101101111100010000;
   assign mem[15766] = 32'b00000000001001011001101101101100;
   assign mem[15767] = 32'b11110101101011111101001111010000;
   assign mem[15768] = 32'b11111000101101001000000110101000;
   assign mem[15769] = 32'b00000011000101111111001010111100;
   assign mem[15770] = 32'b00000011001110101000000110000000;
   assign mem[15771] = 32'b00000101000010100111110011100000;
   assign mem[15772] = 32'b00000100010101101100110100111000;
   assign mem[15773] = 32'b11111100000001000101111101000100;
   assign mem[15774] = 32'b00000011011011111110001111101100;
   assign mem[15775] = 32'b11111101111111001110101101110100;
   assign mem[15776] = 32'b11111010111011101000001011110000;
   assign mem[15777] = 32'b11111111011010001010011011111001;
   assign mem[15778] = 32'b11111101111001011101101011111000;
   assign mem[15779] = 32'b11111111110100101110110110010100;
   assign mem[15780] = 32'b11110111000011001110101111010000;
   assign mem[15781] = 32'b00001001011011111111100100110000;
   assign mem[15782] = 32'b00001110111100100101101011110000;
   assign mem[15783] = 32'b11110011000010111000100111110000;
   assign mem[15784] = 32'b00001010101101010010100001110000;
   assign mem[15785] = 32'b11110111011011100010111111110000;
   assign mem[15786] = 32'b11111100101011011110101101100100;
   assign mem[15787] = 32'b11111011110010001101011111000000;
   assign mem[15788] = 32'b11110110010111111101110011110000;
   assign mem[15789] = 32'b11111111111000110010001101000000;
   assign mem[15790] = 32'b11110101111111000001111010010000;
   assign mem[15791] = 32'b00000100000000000001100111010000;
   assign mem[15792] = 32'b11111100011111000111001111000100;
   assign mem[15793] = 32'b00000011011011001010101001001100;
   assign mem[15794] = 32'b00000000000000101000011101011100;
   assign mem[15795] = 32'b00000000011000010111010000100100;
   assign mem[15796] = 32'b00000011010000011001101000101000;
   assign mem[15797] = 32'b11110111100100001001001010000000;
   assign mem[15798] = 32'b00000101100000110111101111100000;
   assign mem[15799] = 32'b11111100111011000100110101111100;
   assign mem[15800] = 32'b11111100111111101100011011000100;
   assign mem[15801] = 32'b00000011101010100011111011101100;
   assign mem[15802] = 32'b00000010100010001101101111001100;
   assign mem[15803] = 32'b11110100101010111101101101000000;
   assign mem[15804] = 32'b00000110111000110111001100000000;
   assign mem[15805] = 32'b11111000011010100000010000101000;
   assign mem[15806] = 32'b11110001111111000001111110100000;
   assign mem[15807] = 32'b00000100010000111011111000010000;
   assign mem[15808] = 32'b11111111100111000100010110011010;
   assign mem[15809] = 32'b00001011110000010010010001000000;
   assign mem[15810] = 32'b11101100011100101110111000100000;
   assign mem[15811] = 32'b00001001010101010100000011010000;
   assign mem[15812] = 32'b00000001101001010101010011011100;
   assign mem[15813] = 32'b00000111001001100001101100110000;
   assign mem[15814] = 32'b11111011110111000111000110001000;
   assign mem[15815] = 32'b11111001001110110010011001100000;
   assign mem[15816] = 32'b00000010011111011101011101001100;
   assign mem[15817] = 32'b11110010010110101011101000010000;
   assign mem[15818] = 32'b00001000111011000000110010110000;
   assign mem[15819] = 32'b11110111000110101000001110110000;
   assign mem[15820] = 32'b11111101011010100110010111001000;
   assign mem[15821] = 32'b00000111001110101100110111110000;
   assign mem[15822] = 32'b00001000101100101001111110110000;
   assign mem[15823] = 32'b11110100001101010101011100100000;
   assign mem[15824] = 32'b00000100010001100110010010011000;
   assign mem[15825] = 32'b00000000011101110000011011101110;
   assign mem[15826] = 32'b11111000001101010110000101100000;
   assign mem[15827] = 32'b11111000001111001011000000011000;
   assign mem[15828] = 32'b11110100110100000101111110010000;
   assign mem[15829] = 32'b00000001101101000100101110010110;
   assign mem[15830] = 32'b00000010110011011110111010100000;
   assign mem[15831] = 32'b11111111100111000001000000011101;
   assign mem[15832] = 32'b11111100111011101000110000011000;
   assign mem[15833] = 32'b11111111101000111001101000101011;
   assign mem[15834] = 32'b11111101110001011011100001000000;
   assign mem[15835] = 32'b00000010011110010100011101110000;
   assign mem[15836] = 32'b00000010110111010111001111000000;
   assign mem[15837] = 32'b00000010110111010111000011010100;
   assign mem[15838] = 32'b11111110011100101101011000011100;
   assign mem[15839] = 32'b00000000011000111010101111101110;
   assign mem[15840] = 32'b00000011101010000011100101101100;
   assign mem[15841] = 32'b00000000110101000110010110011011;
   assign mem[15842] = 32'b00000111101110101011111111111000;
   assign mem[15843] = 32'b00000010001001110111110111010100;
   assign mem[15844] = 32'b00000000101001111010110110110101;
   assign mem[15845] = 32'b11111001001000101001111101101000;
   assign mem[15846] = 32'b11111110101100001101111101111000;
   assign mem[15847] = 32'b00000011000101001011101101000000;
   assign mem[15848] = 32'b11111110111001001010010101101010;
   assign mem[15849] = 32'b11111101111101010101000110010100;
   assign mem[15850] = 32'b00000110001101110010100100000000;
   assign mem[15851] = 32'b11111011010101001101110110100000;
   assign mem[15852] = 32'b00000011111000000000000000101100;
   assign mem[15853] = 32'b00000001000001100010001100110110;
   assign mem[15854] = 32'b11111111010111011011011001110101;
   assign mem[15855] = 32'b00000011010100011010110010111100;
   assign mem[15856] = 32'b11110101001101101011100101110000;
   assign mem[15857] = 32'b11101111101000001011001001100000;
   assign mem[15858] = 32'b00000011101101010110111111111000;
   assign mem[15859] = 32'b11111011000100101000111000100000;
   assign mem[15860] = 32'b11111100101100001101001101101100;
   assign mem[15861] = 32'b11101011010001000001010010100000;
   assign mem[15862] = 32'b11111100111011100000000011110000;
   assign mem[15863] = 32'b00001001010100010010101110010000;
   assign mem[15864] = 32'b11111000100001010101001011010000;
   assign mem[15865] = 32'b00001000010110000100001110110000;
   assign mem[15866] = 32'b00000111101110011010000010011000;
   assign mem[15867] = 32'b11110100011111100100111111110000;
   assign mem[15868] = 32'b00000100010101001001111011100000;
   assign mem[15869] = 32'b11110111101010110111010001100000;
   assign mem[15870] = 32'b11110110001100101110111001010000;
   assign mem[15871] = 32'b00000011111101111000111111010100;
   assign mem[15872] = 32'b00000100010010000110010010100000;
   assign mem[15873] = 32'b11110000110011100111110010010000;
   assign mem[15874] = 32'b11111111011011101000010001001101;
   assign mem[15875] = 32'b00001011100010010100111110000000;
   assign mem[15876] = 32'b11101010101000101100101000000000;
   assign mem[15877] = 32'b11111000100010101100001110111000;
   assign mem[15878] = 32'b11111100000010110010000100011100;
   assign mem[15879] = 32'b00001011101010101001110101110000;
   assign mem[15880] = 32'b11111110010111010100111110111000;
   assign mem[15881] = 32'b00001010101110000001001110000000;
   assign mem[15882] = 32'b00000111000111110000001111101000;
   assign mem[15883] = 32'b11110110000001101010000111010000;
   assign mem[15884] = 32'b00000110011001010000100011100000;
   assign mem[15885] = 32'b11111011001111110011001010110000;
   assign mem[15886] = 32'b00000000000110100111001001000100;
   assign mem[15887] = 32'b11111000010001111100111011100000;
   assign mem[15888] = 32'b00000011100010100001010110101100;
   assign mem[15889] = 32'b00000000101110010110001101111111;
   assign mem[15890] = 32'b00000011011110110010011011111000;
   assign mem[15891] = 32'b00000010011110111010001111010000;
   assign mem[15892] = 32'b00001001000000001011110000100000;
   assign mem[15893] = 32'b11111001110101101010110111100000;
   assign mem[15894] = 32'b00001000010000001110100011100000;
   assign mem[15895] = 32'b11110110110001100010011110010000;
   assign mem[15896] = 32'b00000011010011111101011101010000;
   assign mem[15897] = 32'b11111100011110100100011101000100;
   assign mem[15898] = 32'b00000101100001011000101001000000;
   assign mem[15899] = 32'b11111011001110000101001100110000;
   assign mem[15900] = 32'b00000011010011011011101101000000;
   assign mem[15901] = 32'b00000001011001100000000010011100;
   assign mem[15902] = 32'b00000010001000101111110111010000;
   assign mem[15903] = 32'b11111110010111110111010111100010;
   assign mem[15904] = 32'b11110111110001010101011100110000;
   assign mem[15905] = 32'b11111010101111010001100010011000;
   assign mem[15906] = 32'b11111010001110100000000110100000;
   assign mem[15907] = 32'b11111000010111100101101100101000;
   assign mem[15908] = 32'b00001001111101011000100101010000;
   assign mem[15909] = 32'b11111001101100111100111100011000;
   assign mem[15910] = 32'b11111111011111111001101111111001;
   assign mem[15911] = 32'b11111010110001010111000110011000;
   assign mem[15912] = 32'b11111100111111110011100101001000;
   assign mem[15913] = 32'b00000011000100111100001011111000;
   assign mem[15914] = 32'b11110111101001111001110101110000;
   assign mem[15915] = 32'b00000001011110011101101011110000;
   assign mem[15916] = 32'b00000000110010011001110010010011;
   assign mem[15917] = 32'b11111011100000110111001011110000;
   assign mem[15918] = 32'b00000100111010011100100101011000;
   assign mem[15919] = 32'b11111110001101111001000011110100;
   assign mem[15920] = 32'b11111111011101110001101111000011;
   assign mem[15921] = 32'b00000100000100111100101001001000;
   assign mem[15922] = 32'b11111101001101010010100111111100;
   assign mem[15923] = 32'b11111100101110000011101001101000;
   assign mem[15924] = 32'b11111010101010100101110001100000;
   assign mem[15925] = 32'b00000010011010010001100100010000;
   assign mem[15926] = 32'b00000001011101001000001011000100;
   assign mem[15927] = 32'b11111000000010001000101010000000;
   assign mem[15928] = 32'b00000100101001011100010101101000;
   assign mem[15929] = 32'b11111111000111011011011011000110;
   assign mem[15930] = 32'b11111010110011101011010100010000;
   assign mem[15931] = 32'b00000011001010001101001001110000;
   assign mem[15932] = 32'b00001000100010111011110101000000;
   assign mem[15933] = 32'b11111100000111010011010100100000;
   assign mem[15934] = 32'b00000111100110000110100110100000;
   assign mem[15935] = 32'b11111011110001011001110011000000;
   assign mem[15936] = 32'b11111101111000110000011010111100;
   assign mem[15937] = 32'b11110111110001110010111011010000;
   assign mem[15938] = 32'b11110100101000001101100010000000;
   assign mem[15939] = 32'b11111100101000110111101001001100;
   assign mem[15940] = 32'b11101111001100010100111111000000;
   assign mem[15941] = 32'b00000110000010111011110000001000;
   assign mem[15942] = 32'b00000110001100011101110110111000;
   assign mem[15943] = 32'b00000010010111001000011011110000;
   assign mem[15944] = 32'b11111011010111101100010101001000;
   assign mem[15945] = 32'b11111000001100000110110110000000;
   assign mem[15946] = 32'b11111111001100110111010000011010;
   assign mem[15947] = 32'b11101110111111011100101011000000;
   assign mem[15948] = 32'b00000111001101001001100010001000;
   assign mem[15949] = 32'b00000000110101000111111011100111;
   assign mem[15950] = 32'b11110100110100001001001010010000;
   assign mem[15951] = 32'b11111111110101011001110111111111;
   assign mem[15952] = 32'b00000011110111000011110100001000;
   assign mem[15953] = 32'b00000101101010000010011100011000;
   assign mem[15954] = 32'b11111110100101111101001011110000;
   assign mem[15955] = 32'b00000010100011001110010011100100;
   assign mem[15956] = 32'b00000000010011000100111011011011;
   assign mem[15957] = 32'b11110001110111101101100010000000;
   assign mem[15958] = 32'b00001010101000100101101000100000;
   assign mem[15959] = 32'b11111111011100100110110010010010;
   assign mem[15960] = 32'b00001010100011011010110101010000;
   assign mem[15961] = 32'b11111011111000100100111000111000;
   assign mem[15962] = 32'b00001010001100001000100010110000;
   assign mem[15963] = 32'b11110010001101011010101000010000;
   assign mem[15964] = 32'b00001010100101100110011111010000;
   assign mem[15965] = 32'b11111110101110111110100011110100;
   assign mem[15966] = 32'b00000001111110110001001110111010;
   assign mem[15967] = 32'b11110101111101011111110000010000;
   assign mem[15968] = 32'b11110110111000000000110001000000;
   assign mem[15969] = 32'b11111001000011010000111111000000;
   assign mem[15970] = 32'b00000100101111010101110111111000;
   assign mem[15971] = 32'b11111101100101011010110001100100;
   assign mem[15972] = 32'b00000101010111101110100101101000;
   assign mem[15973] = 32'b00000101001010011100101010000000;
   assign mem[15974] = 32'b11111101010111111010000110000000;
   assign mem[15975] = 32'b00000010110100011001111000101000;
   assign mem[15976] = 32'b11110101110101111101100111010000;
   assign mem[15977] = 32'b11110110110101011110000111110000;
   assign mem[15978] = 32'b11111100010111101111101100010000;
   assign mem[15979] = 32'b11111111110001011000101110101101;
   assign mem[15980] = 32'b11110011111011010000010110000000;
   assign mem[15981] = 32'b00000001110001001101001111001000;
   assign mem[15982] = 32'b11111111100010010001101111100110;
   assign mem[15983] = 32'b11111011101111010100100000000000;
   assign mem[15984] = 32'b00001001001010100011000011000000;
   assign mem[15985] = 32'b00000011011110110001011010110100;
   assign mem[15986] = 32'b11101111010101011110100101100000;
   assign mem[15987] = 32'b11111000010101000011010010000000;
   assign mem[15988] = 32'b11111101110010111000111101000000;
   assign mem[15989] = 32'b00001011101000000101000101110000;
   assign mem[15990] = 32'b11111000010101000010000000000000;
   assign mem[15991] = 32'b11111110110100101100110111111000;
   assign mem[15992] = 32'b11110011000110100110001011000000;
   assign mem[15993] = 32'b11111101001011111010110000001100;
   assign mem[15994] = 32'b11111101110110111111111000010000;
   assign mem[15995] = 32'b00001000000110011000001100010000;
   assign mem[15996] = 32'b11110111101111000100001000100000;
   assign mem[15997] = 32'b11111001101011100100010100010000;
   assign mem[15998] = 32'b00000010101010110010101110010000;
   assign mem[15999] = 32'b11111111101011001100101101000010;


endmodule
