//	5-bit address is expected.
//	Contains 18 numbers (1/1 to 1/18).
//
//	delta = 0.0045 >= 2^-8
//	Therefore, values are provided with 31 fractional bit precision, which is more than enough. 
module ExpTaylorLut
#(parameter
	DATA_WIDTH = 32,
	FRACTION_BITS = 30
)
(
	adr,
	val
);

input	[4:0]					adr;
output	[DATA_WIDTH-1:0]		val;

wire	[31:0]					mem[0:31];
wire	[2*DATA_WIDTH+32-1:0]	intermediate;
wire	[DATA_WIDTH-1:0]		zero;

assign		zero			=	{DATA_WIDTH{1'b0}};
assign		intermediate	=	{zero, mem[adr], zero};
localparam	NEW_FRAC_BITS	=	31 + DATA_WIDTH;
localparam	EXTRA_FRAC_BITS	=	NEW_FRAC_BITS - FRACTION_BITS;
assign		val				=	intermediate[DATA_WIDTH + EXTRA_FRAC_BITS - 1 : EXTRA_FRAC_BITS];

assign	mem[0]	=	32'b0_0000000000000000000000000000000;

assign	mem[1]	=	32'b1_0000000000000000000000000000000;
assign	mem[2]	=	32'b0_1000000000000000000000000000000;
assign	mem[3]	=	32'b0_0101010101010101010101010101010;
assign	mem[4]	=	32'b0_0100000000000000000000000000000;
assign	mem[5]	=	32'b0_0011001100110011001100110011001;
assign	mem[6]	=	32'b0_0010101010101010101010101010101;
assign	mem[7]	=	32'b0_0010010010010010010010010010010;
assign	mem[8]	=	32'b0_0010000000000000000000000000000;
assign	mem[9]	=	32'b0_0001110001110001110001110001110;
assign	mem[10]	=	32'b0_0001100110011001100110011001100;
assign	mem[11]	=	32'b0_0001011101000101110100010111010;
assign	mem[12]	=	32'b0_0001010101010101010101010101010;
assign	mem[13]	=	32'b0_0001001110110001001110110001001;
assign	mem[14]	=	32'b0_0001001001001001001001001001001;
assign	mem[15]	=	32'b0_0001000100010001000100010001000;
assign	mem[16]	=	32'b0_0001000000000000000000000000000;
assign	mem[17]	=	32'b0_0000111100001111000011110000111;
assign	mem[18]	=	32'b0_0000111000111000111000111000111;

assign	mem[19]	=	32'b0_0000000000000000000000000000000;
assign	mem[20]	=	32'b0_0000000000000000000000000000000;
assign	mem[21]	=	32'b0_0000000000000000000000000000000;
assign	mem[22]	=	32'b0_0000000000000000000000000000000;
assign	mem[23]	=	32'b0_0000000000000000000000000000000;
assign	mem[24]	=	32'b0_0000000000000000000000000000000;
assign	mem[25]	=	32'b0_0000000000000000000000000000000;
assign	mem[20]	=	32'b0_0000000000000000000000000000000;
assign	mem[27]	=	32'b0_0000000000000000000000000000000;
assign	mem[28]	=	32'b0_0000000000000000000000000000000;
assign	mem[29]	=	32'b0_0000000000000000000000000000000;
assign	mem[30]	=	32'b0_0000000000000000000000000000000;
assign	mem[31]	=	32'b0_0000000000000000000000000000000;

endmodule