module DenseWeightLut (
    clk,
    adr,
    dataIn,
    dataOut
);

    localparam WORD_SIZE = 32, LENGTH_SIZE = 10;

    localparam ADR_SIZE = $clog2(LENGTH_SIZE);
    input                   clk, wr;
    input   [ADR_SIZE-1:0]  adr;
    input   [WORD_SIZE-1:0] dataIn;
    output  [WORD_SIZE-1:0] dataOut;

    wire [WORD_SIZE-1:0] mem [0:LENGTH_SIZE-1];

    assign dataOut = mem[adr];

   assign mem[31:0] = 32'b11110011001111111111011101000000;
   assign mem[63:32] = 32'b11111010000001101111101000101000;
   assign mem[95:64] = 32'b00000010001111010010011101111100;
   assign mem[127:96] = 32'b00001101010100001111111011110000;
   assign mem[159:128] = 32'b00000111010101011001101000010000;
   assign mem[191:160] = 32'b11110100011101011101011011000000;
   assign mem[223:192] = 32'b00000010001001101100110010101000;
   assign mem[255:224] = 32'b00000101011110010111100011000000;
   assign mem[287:256] = 32'b11111000011111110001101011000000;
   assign mem[319:288] = 32'b11110001010101100110110000110000;
   assign mem[351:320] = 32'b11111010101110111000000010011000;
   assign mem[383:352] = 32'b00000000011011110110101110100010;
   assign mem[415:384] = 32'b00010000001101101011110110100000;
   assign mem[447:416] = 32'b11111000001111011111110110111000;
   assign mem[479:448] = 32'b00000010011011000111011010100000;
   assign mem[511:480] = 32'b11111111000000001111011001101000;
   assign mem[543:512] = 32'b00001011111001010000000101110000;
   assign mem[575:544] = 32'b11111101011011110010010100111000;
   assign mem[607:576] = 32'b11110010110000110000011001010000;
   assign mem[639:608] = 32'b11110110110000010100110111010000;
   assign mem[671:640] = 32'b11111101011100101110001011010000;
   assign mem[703:672] = 32'b00001010110000001000110001010000;
   assign mem[735:704] = 32'b11110110011000001111010001110000;
   assign mem[767:736] = 32'b00000101100000101010011111100000;
   assign mem[799:768] = 32'b00000111011101001000101101010000;
   assign mem[831:800] = 32'b11111110110001110000000111000100;
   assign mem[863:832] = 32'b00000000110001110101001110001100;
   assign mem[895:864] = 32'b00000000101010010101010001000100;
   assign mem[927:896] = 32'b11111110000000111001110001001010;
   assign mem[959:928] = 32'b11110101101011000100110111100000;
   assign mem[991:960] = 32'b00000010011110101111011110111100;
   assign mem[1023:992] = 32'b00000011111001100010001001000100;
   assign mem[1055:1024] = 32'b00001000111100011101110000110000;
   assign mem[1087:1056] = 32'b00000100001001100100010011001000;
   assign mem[1119:1088] = 32'b11111010101101011101101111010000;
   assign mem[1151:1120] = 32'b11111000010101010011001110101000;
   assign mem[1183:1152] = 32'b11111001100001100111111001000000;
   assign mem[1215:1184] = 32'b11111000010001100001001101111000;
   assign mem[1247:1216] = 32'b11110110010011110110100000110000;
   assign mem[1279:1248] = 32'b11111001100101100010011111101000;
   assign mem[1311:1280] = 32'b00000001010100111100111010000000;
   assign mem[1343:1312] = 32'b00000001100010110001111110011100;
   assign mem[1375:1344] = 32'b11111011000000011001000011000000;
   assign mem[1407:1376] = 32'b00000011000000001010010011000000;
   assign mem[1439:1408] = 32'b11111101001011111101011110110100;
   assign mem[1471:1440] = 32'b11111001001111010110100100110000;
   assign mem[1503:1472] = 32'b11111010110100001110001001110000;
   assign mem[1535:1504] = 32'b11111011110001101011101100101000;
   assign mem[1567:1536] = 32'b00000011000001110110101101100100;
   assign mem[1599:1568] = 32'b00000001100000000011111101000110;
   assign mem[1631:1600] = 32'b11111000110100011111010101100000;
   assign mem[1663:1632] = 32'b11111110001110011111001101100000;
   assign mem[1695:1664] = 32'b11110111011001010111100011110000;
   assign mem[1727:1696] = 32'b00000001010110101100111100110110;
   assign mem[1759:1728] = 32'b11111001011000100110101100110000;
   assign mem[1791:1760] = 32'b11111110100011011111011111001000;
   assign mem[1823:1792] = 32'b00000000011010011110111110110101;
   assign mem[1855:1824] = 32'b00000011100100001010101011011100;
   assign mem[1887:1856] = 32'b00001001111100101001001010010000;
   assign mem[1919:1888] = 32'b11111001111100110011011010010000;
   assign mem[1951:1920] = 32'b00000000100010111010110100110000;
   assign mem[1983:1952] = 32'b11111111001001000010110110000111;
   assign mem[2015:1984] = 32'b11111110101110001101100101010100;
   assign mem[2047:2016] = 32'b11111100101011000110100110111000;
   assign mem[2079:2048] = 32'b00000011001000110101000101000000;
   assign mem[2111:2080] = 32'b00000101010000010111010111011000;
   assign mem[2143:2112] = 32'b00000011001101001101101101010100;
   assign mem[2175:2144] = 32'b00000011011000111001000110100000;
   assign mem[2207:2176] = 32'b00000101001101111010101100000000;
   assign mem[2239:2208] = 32'b11111011111101110101001100101000;
   assign mem[2271:2240] = 32'b11111111111010111001001010100000;
   assign mem[2303:2272] = 32'b11111001101100101000001000110000;
   assign mem[2335:2304] = 32'b11111110111011111110011011011000;
   assign mem[2367:2336] = 32'b00000011111011111101111101000100;
   assign mem[2399:2368] = 32'b11111100111011111010101000000000;
   assign mem[2431:2400] = 32'b00000010001100101011110010000100;
   assign mem[2463:2432] = 32'b00000011111000101011110100000100;
   assign mem[2495:2464] = 32'b11111011101000101111111111111000;
   assign mem[2527:2496] = 32'b11110110110010100110110010100000;
   assign mem[2559:2528] = 32'b11111010111010010101011010001000;
   assign mem[2591:2560] = 32'b00000011110110000001011010110100;
   assign mem[2623:2592] = 32'b00001001000010111011010000010000;
   assign mem[2655:2624] = 32'b11111100110110010100011011000000;
   assign mem[2687:2656] = 32'b00000001101101011000001111110010;
   assign mem[2719:2688] = 32'b00000011111011111111010100010000;
   assign mem[2751:2720] = 32'b11111101100001010100000111010000;
   assign mem[2783:2752] = 32'b11111001001100000001100101100000;
   assign mem[2815:2784] = 32'b00000110001100010011010101001000;
   assign mem[2847:2816] = 32'b00000001111000011101001110101010;
   assign mem[2879:2848] = 32'b00000001011110100011111011011100;
   assign mem[2911:2880] = 32'b00000001010111100010110011000000;
   assign mem[2943:2912] = 32'b11111001101011100010111000000000;
   assign mem[2975:2944] = 32'b11111101110000110101010011010000;
   assign mem[3007:2976] = 32'b11111010001000001110110010100000;
   assign mem[3039:3008] = 32'b11111100110111101011100010010000;
   assign mem[3071:3040] = 32'b11111100000010000010111001011100;
   assign mem[3103:3072] = 32'b00000111101000100111100000110000;
   assign mem[3135:3104] = 32'b11111110100011000010110100000100;
   assign mem[3167:3136] = 32'b00000001000001111011100101111110;
   assign mem[3199:3168] = 32'b00000000101010110011110111000010;
   assign mem[3231:3200] = 32'b11111111101011111011001110011101;
   assign mem[3263:3232] = 32'b11111100011101101011011000000000;
   assign mem[3295:3264] = 32'b00000101101100000100010011110000;
   assign mem[3327:3296] = 32'b00000011111100010111110111011000;
   assign mem[3359:3328] = 32'b11111001101101110110001110010000;
   assign mem[3391:3360] = 32'b11111011101000111001111010101000;
   assign mem[3423:3392] = 32'b00001000110100111001100011100000;
   assign mem[3455:3424] = 32'b11111100110010001000011000111100;
   assign mem[3487:3456] = 32'b11111101001001001111101101111000;
   assign mem[3519:3488] = 32'b11111110011111000100111011101110;
   assign mem[3551:3520] = 32'b11110110100011011000101100110000;
   assign mem[3583:3552] = 32'b00000010101011100010100010110100;
   assign mem[3615:3584] = 32'b11111100000010100110100100101000;
   assign mem[3647:3616] = 32'b00000100100110001010010101001000;
   assign mem[3679:3648] = 32'b00000010111111001011101111100100;
   assign mem[3711:3680] = 32'b00000001010111101011000101010000;
   assign mem[3743:3712] = 32'b11111110111101111110001100000000;
   assign mem[3775:3744] = 32'b00000111101111101100011001000000;
   assign mem[3807:3776] = 32'b11111100000100100011110110100000;
   assign mem[3839:3808] = 32'b11110100001011011101110100110000;
   assign mem[3871:3840] = 32'b11111111000100001111010010001111;
   assign mem[3903:3872] = 32'b11111010010101110001001101011000;
   assign mem[3935:3904] = 32'b00000001010000100110111110011100;
   assign mem[3967:3936] = 32'b00000100001010101011000111100000;
   assign mem[3999:3968] = 32'b11111101000101000100101011111100;
   assign mem[4031:4000] = 32'b11111101000000011110011000011000;
   assign mem[4063:4032] = 32'b11110101101100110010000101100000;
   assign mem[4095:4064] = 32'b00000100010000110000001001110000;
   assign mem[4127:4096] = 32'b11111100001001111111111010111000;
   assign mem[4159:4128] = 32'b11111100111100011000000100100100;
   assign mem[4191:4160] = 32'b00000011100111110001010111011000;
   assign mem[4223:4192] = 32'b00001100110100010101100110110000;
   assign mem[4255:4224] = 32'b11110111111000111101011010110000;
   assign mem[4287:4256] = 32'b00000011000100010001110001100100;
   assign mem[4319:4288] = 32'b11111111111111010101000000000001;
   assign mem[4351:4320] = 32'b11111011000011101000001001010000;
   assign mem[4383:4352] = 32'b11110001111100110100100001010000;
   assign mem[4415:4384] = 32'b00000100000111111111011100111000;
   assign mem[4447:4416] = 32'b11111111110001011101110010101100;
   assign mem[4479:4448] = 32'b00000001110011010110000111101000;
   assign mem[4511:4480] = 32'b00000001000001010110101010111110;
   assign mem[4543:4512] = 32'b11111110110001001001111000001000;
   assign mem[4575:4544] = 32'b00000000100000010001101010011100;
   assign mem[4607:4576] = 32'b00000110110101101100101000010000;
   assign mem[4639:4608] = 32'b00000110010111000101101011101000;
   assign mem[4671:4640] = 32'b11110111010110011100111100110000;
   assign mem[4703:4672] = 32'b11111011111010011101000001001000;
   assign mem[4735:4704] = 32'b00000000110011101110000101001010;
   assign mem[4767:4736] = 32'b11111110110100011000000001111010;
   assign mem[4799:4768] = 32'b11111001111100011011110001011000;
   assign mem[4831:4800] = 32'b00000010100000100000001011100100;
   assign mem[4863:4832] = 32'b11111011000101001100011100110000;
   assign mem[4895:4864] = 32'b00000000101011011100110101011011;
   assign mem[4927:4896] = 32'b00000010001001100001110111011100;
   assign mem[4959:4928] = 32'b11111011011100000011100000010000;
   assign mem[4991:4960] = 32'b11111100100100100010010101111000;
   assign mem[5023:4992] = 32'b00000101111100001100010110111000;
   assign mem[5055:5024] = 32'b11110111111111011011110010100000;
   assign mem[5087:5056] = 32'b00000101000010110001111100010000;
   assign mem[5119:5088] = 32'b00000001111110111011101111111100;
   assign mem[5151:5120] = 32'b11110111001011111100101010000000;
   assign mem[5183:5152] = 32'b00000001010100011010110001011010;
   assign mem[5215:5184] = 32'b00001011011100010111100101000000;
   assign mem[5247:5216] = 32'b00000010010111101110011101101000;
   assign mem[5279:5248] = 32'b11111011101111010101100100111000;
   assign mem[5311:5280] = 32'b11101011010011001001111001100000;
   assign mem[5343:5312] = 32'b00000010110100100011111110000100;
   assign mem[5375:5344] = 32'b00000100011000011010111001001000;
   assign mem[5407:5376] = 32'b11110100111101010010110101110000;
   assign mem[5439:5408] = 32'b11110011010000111100001011100000;
   assign mem[5471:5440] = 32'b11111110101110011111101101000100;
   assign mem[5503:5472] = 32'b00000111100000001101100010011000;
   assign mem[5535:5504] = 32'b11111001001010001111111101001000;
   assign mem[5567:5536] = 32'b00000101011111110010011011010000;
   assign mem[5599:5568] = 32'b00000000100001010111001110100111;
   assign mem[5631:5600] = 32'b11111111011111110010110111000111;
   assign mem[5663:5632] = 32'b00000010010100100110101001011000;
   assign mem[5695:5664] = 32'b11111101100000011000010011011100;
   assign mem[5727:5696] = 32'b11111111101011100010001100011011;
   assign mem[5759:5728] = 32'b11110101001011101011111010010000;
   assign mem[5791:5760] = 32'b11111011010111011001010011001000;
   assign mem[5823:5792] = 32'b00000011100000000100100100101000;
   assign mem[5855:5824] = 32'b11111101110001100001101111110100;
   assign mem[5887:5856] = 32'b11111001101110000001000011101000;
   assign mem[5919:5888] = 32'b00001110100111100110110010010000;
   assign mem[5951:5920] = 32'b11110111100000000011011111100000;
   assign mem[5983:5952] = 32'b00000011111111010011110000100100;
   assign mem[6015:5984] = 32'b00000101001000011100010011110000;
   assign mem[6047:6016] = 32'b11101101101010101111001110100000;
   assign mem[6079:6048] = 32'b11101000011011001000110100000000;
   assign mem[6111:6080] = 32'b11111001011100100010111001111000;
   assign mem[6143:6112] = 32'b11111110000111010000111100001110;
   assign mem[6175:6144] = 32'b11111111011011011001110111000111;
   assign mem[6207:6176] = 32'b00000101000010001110100101111000;
   assign mem[6239:6208] = 32'b00001000100000011001011010110000;
   assign mem[6271:6240] = 32'b11111000110111010100111111000000;
   assign mem[6303:6272] = 32'b00000000111011011111110100011110;
   assign mem[6335:6304] = 32'b11110101100111110110010100110000;
   assign mem[6367:6336] = 32'b00000110011100000001011111001000;
   assign mem[6399:6368] = 32'b11111111010110110010010110000111;
   assign mem[6431:6400] = 32'b00000011001011110000110101101100;
   assign mem[6463:6432] = 32'b11111010100010101101101111101000;
   assign mem[6495:6464] = 32'b11111001111101110101011000110000;
   assign mem[6527:6496] = 32'b00000001010110001111110011111010;
   assign mem[6559:6528] = 32'b11111110110001011011010010001000;
   assign mem[6591:6560] = 32'b00000000000010101000011010000111;
   assign mem[6623:6592] = 32'b00001110010010101011000111010000;
   assign mem[6655:6624] = 32'b11110111101110010111101001100000;
   assign mem[6687:6656] = 32'b11111111110101100101110001010101;
   assign mem[6719:6688] = 32'b00000000111001111000000000111011;
   assign mem[6751:6720] = 32'b00000100001111001010000110001000;
   assign mem[6783:6752] = 32'b11111110101101111100010000010110;
   assign mem[6815:6784] = 32'b11111100111110000111011000101100;
   assign mem[6847:6816] = 32'b00000100110011000100000110110000;
   assign mem[6879:6848] = 32'b00000001110011001001011111011010;
   assign mem[6911:6880] = 32'b11110110011101100100011010100000;
   assign mem[6943:6912] = 32'b11111111101110001111100011010110;
   assign mem[6975:6944] = 32'b00000001100011100100111010010000;
   assign mem[7007:6976] = 32'b00000000110110101010010101011111;
   assign mem[7039:7008] = 32'b00000001111101010000101011111000;
   assign mem[7071:7040] = 32'b11110101110000111101000101010000;
   assign mem[7103:7072] = 32'b11111101110101000001100001101000;
   assign mem[7135:7104] = 32'b11111010001010101100111111000000;
   assign mem[7167:7136] = 32'b00000101010001100001001100101000;
   assign mem[7199:7168] = 32'b11111111100110100011110100010011;
   assign mem[7231:7200] = 32'b11111100001111101100100001011000;
   assign mem[7263:7232] = 32'b00001100001100101111011001110000;
   assign mem[7295:7264] = 32'b11110111000001100001110110100000;
   assign mem[7327:7296] = 32'b00000000100100101100011101000101;
   assign mem[7359:7328] = 32'b11110101101100010010110011100000;
   assign mem[7391:7360] = 32'b11111111000101000100010101111100;
   assign mem[7423:7392] = 32'b00001011100000110110111011100000;
   assign mem[7455:7424] = 32'b11110101111011100001001011100000;
   assign mem[7487:7456] = 32'b00000011001101010111100100010100;
   assign mem[7519:7488] = 32'b11111111100011011001101101100100;
   assign mem[7551:7520] = 32'b00000001011101110001000111111010;
   assign mem[7583:7552] = 32'b00001000101001000101010100010000;
   assign mem[7615:7584] = 32'b00000101000001010000101001111000;
   assign mem[7647:7616] = 32'b00000000000100001100111101111001;
   assign mem[7679:7648] = 32'b11110110101011100110010000010000;
   assign mem[7711:7680] = 32'b11111011000001011101100001000000;
   assign mem[7743:7712] = 32'b00001000111101100101000011110000;
   assign mem[7775:7744] = 32'b11110011000010010111101001000000;
   assign mem[7807:7776] = 32'b00000101010010000101111111011000;
   assign mem[7839:7808] = 32'b00000010100010110011110100111100;
   assign mem[7871:7840] = 32'b00000111001010000111101001011000;
   assign mem[7903:7872] = 32'b00000101111001100111011100101000;
   assign mem[7935:7904] = 32'b00000010110010110101111101000000;
   assign mem[7967:7936] = 32'b11111001011101010110101011100000;
   assign mem[7999:7968] = 32'b11110010111101010100110010010000;
   assign mem[8031:8000] = 32'b11111010011110010100101100000000;
   assign mem[8063:8032] = 32'b11111011101000111101010111101000;
   assign mem[8095:8064] = 32'b11111100001001111011000110011100;
   assign mem[8127:8096] = 32'b11111110101011010001010011001100;
   assign mem[8159:8128] = 32'b11111101001001100101001000001100;
   assign mem[8191:8160] = 32'b00000000101110100110111110010111;
   assign mem[8223:8192] = 32'b00001011110000111110000011110000;
   assign mem[8255:8224] = 32'b00000001100101100110001000010000;
   assign mem[8287:8256] = 32'b11111111001011011000110110011110;
   assign mem[8319:8288] = 32'b11111110101110100111101100011100;
   assign mem[8351:8320] = 32'b11101111011101111010101010100000;
   assign mem[8383:8352] = 32'b00000000110100110110100111111110;
   assign mem[8415:8384] = 32'b11111110101011111100011001111000;
   assign mem[8447:8416] = 32'b11110011001110100110110111110000;
   assign mem[8479:8448] = 32'b00000010101001001001010111011000;
   assign mem[8511:8480] = 32'b00000010000011110110011011101100;
   assign mem[8543:8512] = 32'b00001110010100111011111010010000;
   assign mem[8575:8544] = 32'b11110101100000101101010011010000;
   assign mem[8607:8576] = 32'b11111111001100110101011001100001;
   assign mem[8639:8608] = 32'b11101111111111010110010100000000;
   assign mem[8671:8640] = 32'b00000000101110001100011010101101;
   assign mem[8703:8672] = 32'b11111100101001110111000000010100;
   assign mem[8735:8704] = 32'b11111111110000110101000001011101;
   assign mem[8767:8736] = 32'b00000010100100001011010000010000;
   assign mem[8799:8768] = 32'b00000010101110011011110000100100;
   assign mem[8831:8800] = 32'b11111110010100010100111111110100;
   assign mem[8863:8832] = 32'b11111101000001001000011011111100;
   assign mem[8895:8864] = 32'b11111111001110011000101001011011;
   assign mem[8927:8896] = 32'b00000100110000100010111011000000;
   assign mem[8959:8928] = 32'b00000000100111010100101011100111;
   assign mem[8991:8960] = 32'b11111111110011001011101100000001;
   assign mem[9023:8992] = 32'b11111011100100001111100000111000;
   assign mem[9055:9024] = 32'b00000100110111001010111100001000;
   assign mem[9087:9056] = 32'b00001000100110100100100110110000;
   assign mem[9119:9088] = 32'b11111110111100010010000001000000;
   assign mem[9151:9120] = 32'b11111110101110100101001011010010;
   assign mem[9183:9152] = 32'b00000001100001110001010000101000;
   assign mem[9215:9184] = 32'b11111011011010100100110101100000;
   assign mem[9247:9216] = 32'b11111110001110010101110000101100;
   assign mem[9279:9248] = 32'b11111101001111000000111001010100;
   assign mem[9311:9280] = 32'b00000001011011010010001101110110;
   assign mem[9343:9312] = 32'b00000101011010110010001110110000;
   assign mem[9375:9344] = 32'b11111110111100011110101001001000;
   assign mem[9407:9376] = 32'b00000001100001101011010011111000;
   assign mem[9439:9408] = 32'b00000000011100001010011111110110;
   assign mem[9471:9440] = 32'b11111010001100110101011001011000;
   assign mem[9503:9472] = 32'b11111010100110001000000111110000;
   assign mem[9535:9504] = 32'b00000010001110001010100011010100;
   assign mem[9567:9536] = 32'b11111111110110110100010001100001;
   assign mem[9599:9568] = 32'b11111110110010011110010001010000;
   assign mem[9631:9600] = 32'b00000001000111110010100101111110;
   assign mem[9663:9632] = 32'b00000001011011011110010010101000;
   assign mem[9695:9664] = 32'b11111101101110111010110001001000;
   assign mem[9727:9696] = 32'b11110111001100010010111111010000;
   assign mem[9759:9728] = 32'b11111111110000111011000001110000;
   assign mem[9791:9760] = 32'b11111111011011100001011001111100;
   assign mem[9823:9792] = 32'b00001101011110100000101111110000;
   assign mem[9855:9824] = 32'b00000001001011011000000111010010;
   assign mem[9887:9856] = 32'b11111010100111010111001101100000;
   assign mem[9919:9888] = 32'b11101000100001100110000000100000;
   assign mem[9951:9920] = 32'b11111011110001011111011000101000;
   assign mem[9983:9952] = 32'b11111101010011110111000010111000;
   assign mem[10015:9984] = 32'b00000010000001110001110100100000;
   assign mem[10047:10016] = 32'b00000101100100011100100000111000;
   assign mem[10079:10048] = 32'b11111010110001000001001011100000;
   assign mem[10111:10080] = 32'b11101010101101010101101000100000;
   assign mem[10143:10112] = 32'b00000100101010011010111111101000;
   assign mem[10175:10144] = 32'b00000101011001100100100000111000;
   assign mem[10207:10176] = 32'b11110011000110000000100100100000;
   assign mem[10239:10208] = 32'b11110010111011001010111101000000;
   assign mem[10271:10240] = 32'b00000110001000101011000111011000;
   assign mem[10303:10272] = 32'b11110011001110001100000100110000;
   assign mem[10335:10304] = 32'b00000001010100011111101100101100;
   assign mem[10367:10336] = 32'b00000010000010000110100000010000;
   assign mem[10399:10368] = 32'b00000010010011101011010110100000;
   assign mem[10431:10400] = 32'b11111011111101011100111000110000;
   assign mem[10463:10432] = 32'b00000100001101001100110001101000;
   assign mem[10495:10464] = 32'b11111101011010100111010001100000;
   assign mem[10527:10496] = 32'b00000111001010101000011100100000;
   assign mem[10559:10528] = 32'b11110111011111111000001111000000;
   assign mem[10591:10560] = 32'b11111101010000000101100011001100;
   assign mem[10623:10592] = 32'b11111101010110000101010001001100;
   assign mem[10655:10624] = 32'b11111111111011000000010101110100;
   assign mem[10687:10656] = 32'b00000100010000110001011111100000;
   assign mem[10719:10688] = 32'b00000110000000001001100101001000;
   assign mem[10751:10720] = 32'b11111100100101111100110110101100;
   assign mem[10783:10752] = 32'b00001001110101001100101101100000;
   assign mem[10815:10784] = 32'b11110100000000001100010100110000;
   assign mem[10847:10816] = 32'b00000001101101000000110100100110;
   assign mem[10879:10848] = 32'b11111001111011010000010101111000;
   assign mem[10911:10880] = 32'b11110111100001100100000000110000;
   assign mem[10943:10912] = 32'b11111100000000001111010110101100;
   assign mem[10975:10944] = 32'b00000001011000001010001011111010;
   assign mem[11007:10976] = 32'b00000011011000110000101001001100;
   assign mem[11039:11008] = 32'b11111110110111110011010110010100;
   assign mem[11071:11040] = 32'b11110100110010001111111111110000;
   assign mem[11103:11072] = 32'b00001010110100111100101001000000;
   assign mem[11135:11104] = 32'b00000000111101010011010111001110;
   assign mem[11167:11136] = 32'b11110110100000000001001100010000;
   assign mem[11199:11168] = 32'b11101110001001110001001111000000;
   assign mem[11231:11200] = 32'b00000100001111101001011111100000;
   assign mem[11263:11232] = 32'b11110111101100101011111110100000;
   assign mem[11295:11264] = 32'b11111110101000101011001110101100;
   assign mem[11327:11296] = 32'b11111101110100110111000000100100;
   assign mem[11359:11328] = 32'b11111101111001100000110010100100;
   assign mem[11391:11360] = 32'b00000000001100101111000001001010;
   assign mem[11423:11392] = 32'b11111001110111100111011100101000;
   assign mem[11455:11424] = 32'b00000000000010010110011010110011;
   assign mem[11487:11456] = 32'b00001001010010110100111000010000;
   assign mem[11519:11488] = 32'b00000010101010011010110011111000;
   assign mem[11551:11520] = 32'b00000000011000100101010101101101;
   assign mem[11583:11552] = 32'b00000110111011010010101011110000;
   assign mem[11615:11584] = 32'b11111111110111110111111101101101;
   assign mem[11647:11616] = 32'b11111011010101010110110111110000;
   assign mem[11679:11648] = 32'b00000010111000011110110100101100;
   assign mem[11711:11680] = 32'b11111111111000011110000110001100;
   assign mem[11743:11712] = 32'b11110110111101101110100100100000;
   assign mem[11775:11744] = 32'b00000100011000101110100101000000;
   assign mem[11807:11776] = 32'b11111101110111010111000001100100;
   assign mem[11839:11808] = 32'b11111100111001100101110000011100;
   assign mem[11871:11840] = 32'b11111010000110011011110110111000;
   assign mem[11903:11872] = 32'b00001100010111101100101111000000;
   assign mem[11935:11904] = 32'b11110111100101000010000110010000;
   assign mem[11967:11936] = 32'b00001001000000010111101010000000;
   assign mem[11999:11968] = 32'b00000001001010101101010110011100;
   assign mem[12031:12000] = 32'b11111101111010100001100010101000;
   assign mem[12063:12032] = 32'b00000011011001110100001111101100;
   assign mem[12095:12064] = 32'b00001010011001000011001001100000;
   assign mem[12127:12096] = 32'b11111110011001000001111011100110;
   assign mem[12159:12128] = 32'b11110101000110101101001111010000;
   assign mem[12191:12160] = 32'b00000001011011111110111110100000;
   assign mem[12223:12192] = 32'b11111111111001010011010111000000;
   assign mem[12255:12224] = 32'b00000000100000011000111100011100;
   assign mem[12287:12256] = 32'b00000111011111110110101111010000;
   assign mem[12319:12288] = 32'b11111010000110111010001101110000;
   assign mem[12351:12320] = 32'b11111011000000111110101001000000;
   assign mem[12383:12352] = 32'b00000000110101101000110000101110;
   assign mem[12415:12384] = 32'b00000101111111011110101001111000;
   assign mem[12447:12416] = 32'b11110111011101100001010111100000;
   assign mem[12479:12448] = 32'b11111110111110101110101010011100;
   assign mem[12511:12480] = 32'b00000111001011100101110010111000;
   assign mem[12543:12512] = 32'b11111010010110111010001111001000;
   assign mem[12575:12544] = 32'b11111101011010110010101000111000;
   assign mem[12607:12576] = 32'b00000000100110100011001011000110;
   assign mem[12639:12608] = 32'b11111100101011110010010010101100;
   assign mem[12671:12640] = 32'b11111110100111100111011101011010;
   assign mem[12703:12672] = 32'b11111000000001001111110001010000;
   assign mem[12735:12704] = 32'b11111100110010110000001110010100;
   assign mem[12767:12736] = 32'b11111101000100100010001110011000;
   assign mem[12799:12768] = 32'b00000001111110111110011110101000;
   assign mem[12831:12800] = 32'b11111100011111001010001100010000;
   assign mem[12863:12832] = 32'b00001001110011010111101101010000;
   assign mem[12895:12864] = 32'b11111100011001001001101110101100;
   assign mem[12927:12896] = 32'b00000001111001000000001011011100;
   assign mem[12959:12928] = 32'b00000011110001110100110111000100;
   assign mem[12991:12960] = 32'b11111000011110101000110010111000;
   assign mem[13023:12992] = 32'b11111001000111111001000001110000;
   assign mem[13055:13024] = 32'b11111110110110000011110011010100;
   assign mem[13087:13056] = 32'b11111010110010000111100100011000;
   assign mem[13119:13088] = 32'b11110101000101100100011101010000;
   assign mem[13151:13120] = 32'b11110110111000001000111001110000;
   assign mem[13183:13152] = 32'b11111100001000110110100011110100;
   assign mem[13215:13184] = 32'b00000010110111001110000011101000;
   assign mem[13247:13216] = 32'b00000101011101001001010010111000;
   assign mem[13279:13248] = 32'b11110111110011011111101100100000;
   assign mem[13311:13280] = 32'b11110010000010100011001110100000;
   assign mem[13343:13312] = 32'b11111011000000110001110011001000;
   assign mem[13375:13344] = 32'b11111001001011111000010101010000;
   assign mem[13407:13376] = 32'b11111001010100111011101001100000;
   assign mem[13439:13408] = 32'b00000000111010100001011110111011;
   assign mem[13471:13440] = 32'b11111001111100010100110101011000;
   assign mem[13503:13472] = 32'b00000011010101001011100101000100;
   assign mem[13535:13504] = 32'b00000001100111101010001110000110;
   assign mem[13567:13536] = 32'b00000101100110110000101010010000;
   assign mem[13599:13568] = 32'b11111101100010011010000101010000;
   assign mem[13631:13600] = 32'b11101111001010010001010101100000;
   assign mem[13663:13632] = 32'b00000010010100110000101011011100;
   assign mem[13695:13664] = 32'b00000101010000011000101000000000;
   assign mem[13727:13696] = 32'b00000010110110111000011100010100;
   assign mem[13759:13728] = 32'b11111100100110010001010100100000;
   assign mem[13791:13760] = 32'b11110100111100110010101011110000;
   assign mem[13823:13792] = 32'b00000001100100001010011100111110;
   assign mem[13855:13824] = 32'b00000000101011101110110111111000;
   assign mem[13887:13856] = 32'b11111001101001110110001000100000;
   assign mem[13919:13888] = 32'b11111110101011101001111011011010;
   assign mem[13951:13920] = 32'b11111110011010010101011111101000;
   assign mem[13983:13952] = 32'b00010001100001011001101001000000;
   assign mem[14015:13984] = 32'b11111101010000000000110000010000;
   assign mem[14047:14016] = 32'b11111110001000010001100100011000;
   assign mem[14079:14048] = 32'b11111110010111100001100100101000;
   assign mem[14111:14080] = 32'b00000001000000111000000001110100;
   assign mem[14143:14112] = 32'b00000011010100000100011001010000;
   assign mem[14175:14144] = 32'b11111111101000001101110110000000;
   assign mem[14207:14176] = 32'b00000110010100010000101000011000;
   assign mem[14239:14208] = 32'b11111000010100000001110010011000;
   assign mem[14271:14240] = 32'b11111010000100000100101110111000;
   assign mem[14303:14272] = 32'b11111110011001110110111010001000;
   assign mem[14335:14304] = 32'b00000000101110010011111101001011;
   assign mem[14367:14336] = 32'b11111100101100000010100111000100;
   assign mem[14399:14368] = 32'b11111101101101101000111011000100;
   assign mem[14431:14400] = 32'b00000100010011011010000001101000;
   assign mem[14463:14432] = 32'b11111100100100010100111011111000;
   assign mem[14495:14464] = 32'b11111100011000010110000101001100;
   assign mem[14527:14496] = 32'b11111111100110000010001110011010;
   assign mem[14559:14528] = 32'b00000100010000000100001001101000;
   assign mem[14591:14560] = 32'b11111111111011111100000100100100;
   assign mem[14623:14592] = 32'b00000001000100010010110111101110;
   assign mem[14655:14624] = 32'b00000101101100001110010011001000;
   assign mem[14687:14656] = 32'b11111111101000101011000110111110;
   assign mem[14719:14688] = 32'b11111011011011001110001011011000;
   assign mem[14751:14720] = 32'b11111110000100010100001011110000;
   assign mem[14783:14752] = 32'b11110100001110100011100101000000;
   assign mem[14815:14784] = 32'b00000001100000001110001100100110;
   assign mem[14847:14816] = 32'b11111000010111110010010010110000;
   assign mem[14879:14848] = 32'b11111111110101111110010101110111;
   assign mem[14911:14880] = 32'b00000011101010001011111101111000;
   assign mem[14943:14912] = 32'b00001011110000010000111000010000;
   assign mem[14975:14944] = 32'b11111100011110111100011001010100;
   assign mem[15007:14976] = 32'b00000000110011111000100100110111;
   assign mem[15039:15008] = 32'b00000000011001011011010000101101;
   assign mem[15071:15040] = 32'b00000000100101011101010111010011;
   assign mem[15103:15072] = 32'b00000000111100011101011000001000;
   assign mem[15135:15104] = 32'b00000001101100000011011111110110;
   assign mem[15167:15136] = 32'b11111101101111001011010111000000;
   assign mem[15199:15168] = 32'b11111100111100101010111101011000;
   assign mem[15231:15200] = 32'b11111011101111101001111110111000;
   assign mem[15263:15232] = 32'b00000010100111010011010011111100;
   assign mem[15295:15264] = 32'b11111101110000000010101000000100;
   assign mem[15327:15296] = 32'b11111111101011010101010100000100;
   assign mem[15359:15328] = 32'b11111100111110110010000101011100;
   assign mem[15391:15360] = 32'b11111100110111000011101100110000;
   assign mem[15423:15392] = 32'b11111100010111110100000000010000;
   assign mem[15455:15424] = 32'b00000001110101000111100100111010;
   assign mem[15487:15456] = 32'b00000100010110100110110001010000;
   assign mem[15519:15488] = 32'b11111110000101010111100101101100;
   assign mem[15551:15520] = 32'b11111010111110011000110111000000;
   assign mem[15583:15552] = 32'b00000001011111000100101001010110;
   assign mem[15615:15584] = 32'b11111110110101100011110100111100;
   assign mem[15647:15616] = 32'b11111011011101111000011111000000;
   assign mem[15679:15648] = 32'b11111101111001100100100011001100;
   assign mem[15711:15680] = 32'b00000000001000011000111001100101;
   assign mem[15743:15712] = 32'b11110111110010011111001111110000;
   assign mem[15775:15744] = 32'b11111111000110111010011001000100;
   assign mem[15807:15776] = 32'b00000011001011011001101110100100;
   assign mem[15839:15808] = 32'b11111011011010001111100101100000;
   assign mem[15871:15840] = 32'b11111111100100101111101001011010;
   assign mem[15903:15872] = 32'b00001000100001001010001101110000;
   assign mem[15935:15904] = 32'b11111010100010010101001101011000;
   assign mem[15967:15936] = 32'b00000101110011010101000000000000;
   assign mem[15999:15968] = 32'b11111010010100000111000100110000;
   assign mem[16031:16000] = 32'b11111010001001011010100100001000;
   assign mem[16063:16032] = 32'b11111000110000101101101100010000;
   assign mem[16095:16064] = 32'b00000011010100100001111010111000;
   assign mem[16127:16096] = 32'b00000110010001100111010011010000;
   assign mem[16159:16128] = 32'b00001001000000001001101101110000;
   assign mem[16191:16160] = 32'b11111010010000100101100011010000;
   assign mem[16223:16192] = 32'b00000010101000111100110001110000;
   assign mem[16255:16224] = 32'b11101111001100001011100100100000;
   assign mem[16287:16256] = 32'b00000010110000001111101001011000;
   assign mem[16319:16288] = 32'b00000000010101011011100000011010;
   assign mem[16351:16320] = 32'b11111110100101001011010000111100;
   assign mem[16383:16352] = 32'b11111010110000010010011001110000;
   assign mem[16415:16384] = 32'b00000001101000001101000010100010;
   assign mem[16447:16416] = 32'b11111011100101101000111001010000;
   assign mem[16479:16448] = 32'b11111011000110010011010011100000;
   assign mem[16511:16480] = 32'b11111011101000111111000110101000;
   assign mem[16543:16512] = 32'b00001000000101100101001000110000;
   assign mem[16575:16544] = 32'b00000011110011010001101010100100;
   assign mem[16607:16576] = 32'b00000011000011010111000110011100;
   assign mem[16639:16608] = 32'b11111010101001101100111100010000;
   assign mem[16671:16640] = 32'b11111101110010010000010111101100;
   assign mem[16703:16672] = 32'b00000101001000011101110111100000;
   assign mem[16735:16704] = 32'b00000101100101011101001101111000;
   assign mem[16767:16736] = 32'b00000100000100011011010011100000;
   assign mem[16799:16768] = 32'b11110101000110100101011110100000;
   assign mem[16831:16800] = 32'b11101111011000100100111010000000;
   assign mem[16863:16832] = 32'b00000110010101111111101101101000;
   assign mem[16895:16864] = 32'b00000011111110111000011110001000;
   assign mem[16927:16896] = 32'b11110110001100010111111111000000;
   assign mem[16959:16928] = 32'b11110010001011110010110011010000;
   assign mem[16991:16960] = 32'b11111100100101011100011111010100;
   assign mem[17023:16992] = 32'b11111000011010100100010110100000;
   assign mem[17055:17024] = 32'b00000011100100000000101100011100;
   assign mem[17087:17056] = 32'b00000000111001110111100111010011;
   assign mem[17119:17088] = 32'b11111011110000101011101011101000;
   assign mem[17151:17120] = 32'b11110111100001110001100000000000;
   assign mem[17183:17152] = 32'b00000000101100111010001110000001;
   assign mem[17215:17184] = 32'b00000010000111001111001100000000;
   assign mem[17247:17216] = 32'b00000000001111111001100000011001;
   assign mem[17279:17248] = 32'b00000010011100010000110110111100;
   assign mem[17311:17280] = 32'b11111111001011001101010110110000;
   assign mem[17343:17312] = 32'b00000001010010000100110111100110;
   assign mem[17375:17344] = 32'b00000100110010111011101010011000;
   assign mem[17407:17376] = 32'b00000110001111101101100110110000;
   assign mem[17439:17408] = 32'b11110111000010000101011001010000;
   assign mem[17471:17440] = 32'b11101000110011101001110100100000;
   assign mem[17503:17472] = 32'b11111111110001110110111011100111;
   assign mem[17535:17504] = 32'b11111101110110010110011010111000;
   assign mem[17567:17536] = 32'b11110101010101010011111011010000;
   assign mem[17599:17568] = 32'b11110110000100000010000111100000;
   assign mem[17631:17600] = 32'b11111111100111110000100111011000;
   assign mem[17663:17632] = 32'b11111000101010011010110101110000;
   assign mem[17695:17664] = 32'b11111101101101000110010100000000;
   assign mem[17727:17696] = 32'b11111011100110111000110000101000;
   assign mem[17759:17728] = 32'b11111110111110010110101101010100;
   assign mem[17791:17760] = 32'b00000000101001000111100110010100;
   assign mem[17823:17792] = 32'b00000000011011100000110001101110;
   assign mem[17855:17824] = 32'b00000100000100001010111110000000;
   assign mem[17887:17856] = 32'b00001001100000000001101101000000;
   assign mem[17919:17888] = 32'b11111110110110111000010001111000;
   assign mem[17951:17920] = 32'b11111100010000000101111000011000;
   assign mem[17983:17952] = 32'b11111110001111010000100001001000;
   assign mem[18015:17984] = 32'b11111110010100111000000101100100;
   assign mem[18047:18016] = 32'b00000101001001010100111011110000;
   assign mem[18079:18048] = 32'b00000000000101000111000000001011;
   assign mem[18111:18080] = 32'b11111111000010110001010111110110;
   assign mem[18143:18112] = 32'b00000100010111010111000011010000;
   assign mem[18175:18144] = 32'b11111101011001101100101010101000;
   assign mem[18207:18176] = 32'b00000001100000101011010011001100;
   assign mem[18239:18208] = 32'b11111001011001101010100000011000;
   assign mem[18271:18240] = 32'b11111001110001110111100001001000;
   assign mem[18303:18272] = 32'b00001000000010101100111110110000;
   assign mem[18335:18304] = 32'b11111100110011011101011100111000;
   assign mem[18367:18336] = 32'b11111110011110100000111111010110;
   assign mem[18399:18368] = 32'b00000111011010101011110011001000;
   assign mem[18431:18400] = 32'b11111001110110111000001111010000;
   assign mem[18463:18432] = 32'b00000011011010100011000010111000;
   assign mem[18495:18464] = 32'b00000110011111101111110000110000;
   assign mem[18527:18496] = 32'b00000001101010111011101001110110;
   assign mem[18559:18528] = 32'b11101011010100100110100111100000;
   assign mem[18591:18560] = 32'b00000010011111001100111101011100;
   assign mem[18623:18592] = 32'b00000001111111101011100010101110;
   assign mem[18655:18624] = 32'b00000000101010011111110110110011;
   assign mem[18687:18656] = 32'b11111111110101100000011010011000;
   assign mem[18719:18688] = 32'b11111100011010111100011001111000;
   assign mem[18751:18720] = 32'b00000000001010001111111010000011;
   assign mem[18783:18752] = 32'b11110101110101101001010101010000;
   assign mem[18815:18784] = 32'b11111111100100000000010111100101;
   assign mem[18847:18816] = 32'b00000001111011101010010001011010;
   assign mem[18879:18848] = 32'b00000001101011001010111010000000;
   assign mem[18911:18880] = 32'b11111101111000000000111111000000;
   assign mem[18943:18912] = 32'b00000010101001011110110011001000;
   assign mem[18975:18944] = 32'b11111010101100111111011010110000;
   assign mem[19007:18976] = 32'b00000000011110000001000001011110;
   assign mem[19039:19008] = 32'b11111101001000100100010110100000;
   assign mem[19071:19040] = 32'b11111011000011100011101111011000;
   assign mem[19103:19072] = 32'b00000100111110000111100110000000;
   assign mem[19135:19104] = 32'b00000111100110011110000111111000;
   assign mem[19167:19136] = 32'b00000000101110010001100110001110;
   assign mem[19199:19168] = 32'b11111101110011110111110000110100;
   assign mem[19231:19200] = 32'b00000101011000000111010000100000;
   assign mem[19263:19232] = 32'b11111100000000110001001111101000;
   assign mem[19295:19264] = 32'b11111110000110001111011110000100;
   assign mem[19327:19296] = 32'b11111100111110010010100111110100;
   assign mem[19359:19328] = 32'b00000000111110010000011001100111;
   assign mem[19391:19360] = 32'b11111010101110001000111111111000;
   assign mem[19423:19392] = 32'b11111100001110110100110100110000;
   assign mem[19455:19424] = 32'b11111111110110010100110101111000;
   assign mem[19487:19456] = 32'b00000000100110001101111000111111;
   assign mem[19519:19488] = 32'b11111011000010011010100010000000;
   assign mem[19551:19520] = 32'b11111011111110000111101011011000;
   assign mem[19583:19552] = 32'b11111000110010101011111100001000;
   assign mem[19615:19584] = 32'b11111101110101011100100000111000;
   assign mem[19647:19616] = 32'b00000110100011110110000110111000;
   assign mem[19679:19648] = 32'b00000011100100100101100000010100;
   assign mem[19711:19680] = 32'b11111010010001110100101010111000;
   assign mem[19743:19712] = 32'b00000111001001100000010100011000;
   assign mem[19775:19744] = 32'b11111011001111110101001101101000;
   assign mem[19807:19776] = 32'b00000001001100101110110011111000;
   assign mem[19839:19808] = 32'b11111010110011011110001101011000;
   assign mem[19871:19840] = 32'b00000001000111111110100011010110;
   assign mem[19903:19872] = 32'b11111110000101110011001101010110;
   assign mem[19935:19904] = 32'b11111001011000010010001010110000;
   assign mem[19967:19936] = 32'b00000001011011101001111000110010;
   assign mem[19999:19968] = 32'b11111110110001111101111000110000;
   assign mem[20031:20000] = 32'b00000001101001011100111110101110;
   assign mem[20063:20032] = 32'b00000111101100001000101000110000;
   assign mem[20095:20064] = 32'b00000001110110101111101101101010;
   assign mem[20127:20096] = 32'b00000010110000001111010001001100;
   assign mem[20159:20128] = 32'b00000001110001011101011110100010;
   assign mem[20191:20160] = 32'b00000001101010000110100111111100;
   assign mem[20223:20192] = 32'b11111011110100011100100101101000;
   assign mem[20255:20224] = 32'b00000000111101110011100110011010;
   assign mem[20287:20256] = 32'b11111001111101110101111000010000;
   assign mem[20319:20288] = 32'b11111110111100101000111100000100;
   assign mem[20351:20320] = 32'b11111011110101101111110111001000;
   assign mem[20383:20352] = 32'b00000011000011111000100011111100;
   assign mem[20415:20384] = 32'b11110111111100111111111100100000;
   assign mem[20447:20416] = 32'b11111111100110010111000100000111;
   assign mem[20479:20448] = 32'b11111110100010011010101000011010;
   assign mem[20511:20480] = 32'b11111011011110100111101110111000;
   assign mem[20543:20512] = 32'b11111100011011011011010001010000;
   assign mem[20575:20544] = 32'b00000000001010001100010000000101;
   assign mem[20607:20576] = 32'b00000011100110011111000011001000;
   assign mem[20639:20608] = 32'b11111010010000001001011100011000;
   assign mem[20671:20640] = 32'b00001010000111010010000110100000;
   assign mem[20703:20672] = 32'b11101111101100111111000000000000;
   assign mem[20735:20704] = 32'b00000110001011100011001111110000;
   assign mem[20767:20736] = 32'b11111101010000110100101100001100;
   assign mem[20799:20768] = 32'b11111101100101010110111111010000;
   assign mem[20831:20800] = 32'b11111001110000011010011010100000;
   assign mem[20863:20832] = 32'b00000100111111111010000111011000;
   assign mem[20895:20864] = 32'b11111101000001001101101001101100;
   assign mem[20927:20896] = 32'b11111110101111111000011010001000;
   assign mem[20959:20928] = 32'b00001001011011011101010100000000;
   assign mem[20991:20960] = 32'b11110001100001001011101001000000;
   assign mem[21023:20992] = 32'b00000010000100000110101101111000;
   assign mem[21055:21024] = 32'b00001000001111010101100110100000;
   assign mem[21087:21056] = 32'b11111100101001010100100011001000;
   assign mem[21119:21088] = 32'b11101100100111010010001111100000;
   assign mem[21151:21120] = 32'b11111111110110000000100010010001;
   assign mem[21183:21152] = 32'b00001010001010010010110111100000;
   assign mem[21215:21184] = 32'b00001000110100011111010011000000;
   assign mem[21247:21216] = 32'b00000001101100010000001101100010;
   assign mem[21279:21248] = 32'b11111111110000010101111010001010;
   assign mem[21311:21280] = 32'b11111010100011011000001110001000;
   assign mem[21343:21312] = 32'b11110101110001111100010101100000;
   assign mem[21375:21344] = 32'b00000001111111100101001110100000;
   assign mem[21407:21376] = 32'b11111011110000001111111000001000;
   assign mem[21439:21408] = 32'b11110101101110001101010010110000;
   assign mem[21471:21440] = 32'b11110101100100111010111110110000;
   assign mem[21503:21472] = 32'b11111101010011001110011100001000;
   assign mem[21535:21504] = 32'b00000111111010010011100110001000;
   assign mem[21567:21536] = 32'b00000101011110001100100100101000;
   assign mem[21599:21568] = 32'b11111010010111100011001110001000;
   assign mem[21631:21600] = 32'b11100111011011010010010001000000;
   assign mem[21663:21632] = 32'b11110100111110110100001111100000;
   assign mem[21695:21664] = 32'b11111100100111000110001000101100;
   assign mem[21727:21696] = 32'b11111100101110110000001111110000;
   assign mem[21759:21728] = 32'b11111101110011101111001001110000;
   assign mem[21791:21760] = 32'b00000000010111011100011000100100;
   assign mem[21823:21792] = 32'b11111001011111000101110110010000;
   assign mem[21855:21824] = 32'b00001101010110011100010000110000;
   assign mem[21887:21856] = 32'b00000101100001010010010101111000;
   assign mem[21919:21888] = 32'b11111101111010110001010110110100;
   assign mem[21951:21920] = 32'b11110100111011001000100100110000;
   assign mem[21983:21952] = 32'b11111100000000011000100111111000;
   assign mem[22015:21984] = 32'b11110111011000111110100100010000;
   assign mem[22047:22016] = 32'b00000001101010100010010111111110;
   assign mem[22079:22048] = 32'b00000100100000000100100110001000;
   assign mem[22111:22080] = 32'b11111100101011000110101010011100;
   assign mem[22143:22112] = 32'b11111011011110000101010101010000;
   assign mem[22175:22144] = 32'b11111111101100101011011000110011;
   assign mem[22207:22176] = 32'b00001000100100100100111011010000;
   assign mem[22239:22208] = 32'b11110101010010100000100101000000;
   assign mem[22271:22240] = 32'b11111100101101011011101000101000;
   assign mem[22303:22272] = 32'b00001001001110010100100010000000;
   assign mem[22335:22304] = 32'b11111101000100101010001010100100;
   assign mem[22367:22336] = 32'b11111110011001011000011010010010;
   assign mem[22399:22368] = 32'b00000000000011111000011111000100;
   assign mem[22431:22400] = 32'b00000000001111111100110011100000;
   assign mem[22463:22432] = 32'b00000110110100110010100000110000;
   assign mem[22495:22464] = 32'b11111101100111111001101110110100;
   assign mem[22527:22496] = 32'b11110011001001000101110110100000;
   assign mem[22559:22528] = 32'b11111111100010101010111111101111;
   assign mem[22591:22560] = 32'b00000111011010101101100111001000;
   assign mem[22623:22592] = 32'b00001101011101110011110010010000;
   assign mem[22655:22624] = 32'b00000001001100011110010010111100;
   assign mem[22687:22656] = 32'b11111010101110000101000101100000;
   assign mem[22719:22688] = 32'b00000000010010101100000110010010;
   assign mem[22751:22720] = 32'b11110110110111010110001001100000;
   assign mem[22783:22752] = 32'b11111000100101000100001001100000;
   assign mem[22815:22784] = 32'b00000111010000001010001011000000;
   assign mem[22847:22816] = 32'b11111110011111100000101110000000;
   assign mem[22879:22848] = 32'b00000010100111011110011001001100;
   assign mem[22911:22880] = 32'b11111101011100111010110000001000;
   assign mem[22943:22912] = 32'b00001011101010110111100011110000;
   assign mem[22975:22944] = 32'b11110011110011101010101111100000;
   assign mem[23007:22976] = 32'b00000101011100111001001000010000;
   assign mem[23039:23008] = 32'b11111001011010010001111000001000;
   assign mem[23071:23040] = 32'b11111101111100011011000100001100;
   assign mem[23103:23072] = 32'b11111100110110000101000010110000;
   assign mem[23135:23104] = 32'b11111111110110010111011100100000;
   assign mem[23167:23136] = 32'b00000010001110101000111001101000;
   assign mem[23199:23168] = 32'b00000001101000011011111100001110;
   assign mem[23231:23200] = 32'b11111111101011010100111110101001;
   assign mem[23263:23232] = 32'b11110110101010011000110011110000;
   assign mem[23295:23264] = 32'b00000001110001101111011001101110;
   assign mem[23327:23296] = 32'b11111101100111001101101110111100;
   assign mem[23359:23328] = 32'b00000001101100110011011111111000;
   assign mem[23391:23360] = 32'b11111101111111010111100000011100;
   assign mem[23423:23392] = 32'b00000101000110001110011000111000;
   assign mem[23455:23424] = 32'b11111101100100001111110000110100;
   assign mem[23487:23456] = 32'b11111001101111010110001100001000;
   assign mem[23519:23488] = 32'b00000110000001001010110000001000;
   assign mem[23551:23520] = 32'b00000010011110111011100100110000;
   assign mem[23583:23552] = 32'b00000110101000010010010111100000;
   assign mem[23615:23584] = 32'b00000111100111011110000010001000;
   assign mem[23647:23616] = 32'b00000011110111110000010011100000;
   assign mem[23679:23648] = 32'b11111111101110000111111100100101;
   assign mem[23711:23680] = 32'b11111010000101100110100000100000;
   assign mem[23743:23712] = 32'b11110101010010000011010110000000;
   assign mem[23775:23744] = 32'b00000011011101011100111111101000;
   assign mem[23807:23776] = 32'b00000110010000000100000011011000;
   assign mem[23839:23808] = 32'b11110110011010101110011000000000;
   assign mem[23871:23840] = 32'b11111110011100000101111101001000;
   assign mem[23903:23872] = 32'b11110110101011101110000001110000;
   assign mem[23935:23904] = 32'b00000001011001011111101101110100;
   assign mem[23967:23936] = 32'b00000101001101101011011110010000;
   assign mem[23999:23968] = 32'b00001000100001110011101000000000;
   assign mem[24031:24000] = 32'b11110101111100010010001100110000;
   assign mem[24063:24032] = 32'b00001001111001101001100101110000;
   assign mem[24095:24064] = 32'b00000001110010101110010100100100;
   assign mem[24127:24096] = 32'b00000110011100101101010110010000;
   assign mem[24159:24128] = 32'b11111111100101010001011110111111;
   assign mem[24191:24160] = 32'b00000001111101001011101000101000;
   assign mem[24223:24192] = 32'b11110100011000110101001101010000;
   assign mem[24255:24224] = 32'b00001011010000010011000000100000;
   assign mem[24287:24256] = 32'b11111100100000101010001111101100;
   assign mem[24319:24288] = 32'b11100010000110000110100010000000;
   assign mem[24351:24320] = 32'b11111101100111110101101110100100;
   assign mem[24383:24352] = 32'b11110110111010111000010010000000;
   assign mem[24415:24384] = 32'b11111101111100110101100011100100;
   assign mem[24447:24416] = 32'b00000100010110101011101011101000;
   assign mem[24479:24448] = 32'b11111111000110011010011101110101;
   assign mem[24511:24480] = 32'b00000101111111101001010110111000;
   assign mem[24543:24512] = 32'b11101100110011011110100001100000;
   assign mem[24575:24544] = 32'b00000010111011000110110111110000;
   assign mem[24607:24576] = 32'b11111110010000000101101101101000;
   assign mem[24639:24608] = 32'b00000001111100100010101111110100;
   assign mem[24671:24640] = 32'b11111110111011000001010000001000;
   assign mem[24703:24672] = 32'b11111100100010011010101010110000;
   assign mem[24735:24704] = 32'b00000011001010110111010100011000;
   assign mem[24767:24736] = 32'b11111111101010110101011100011011;
   assign mem[24799:24768] = 32'b11111110010010111001001000010100;
   assign mem[24831:24800] = 32'b00000001011001111000101100101000;
   assign mem[24863:24832] = 32'b11110111010110001011101100010000;
   assign mem[24895:24864] = 32'b00000011111111111000100010110100;
   assign mem[24927:24896] = 32'b11111110001101100011000101100100;
   assign mem[24959:24928] = 32'b11111111011101001101001011101011;
   assign mem[24991:24960] = 32'b00000011010001010101001101010000;
   assign mem[25023:24992] = 32'b11111101110011011111111110001000;
   assign mem[25055:25024] = 32'b11111010111101110110000001110000;
   assign mem[25087:25056] = 32'b00000010101001110110110101101000;
   assign mem[25119:25088] = 32'b11110110000011110110101010000000;
   assign mem[25151:25120] = 32'b00000011100010100001110110000000;
   assign mem[25183:25152] = 32'b11111111010001001100100100101001;
   assign mem[25215:25184] = 32'b00000111111001000110011111110000;
   assign mem[25247:25216] = 32'b11111110010101111000110011111000;
   assign mem[25279:25248] = 32'b00000011010110001000010110010100;
   assign mem[25311:25280] = 32'b00000001000010010111011111110000;
   assign mem[25343:25312] = 32'b11111011000100110111011011100000;
   assign mem[25375:25344] = 32'b11111110001100101010110110011110;
   assign mem[25407:25376] = 32'b11111001111110011110001101011000;
   assign mem[25439:25408] = 32'b00000000111110001001011000111110;
   assign mem[25471:25440] = 32'b11111011110010110100100100010000;
   assign mem[25503:25472] = 32'b00000010010100100001111010000100;
   assign mem[25535:25504] = 32'b11111101000001110101111000000000;
   assign mem[25567:25536] = 32'b00000001100100101111111010010100;
   assign mem[25599:25568] = 32'b11111110110110101001011110011010;
   assign mem[25631:25600] = 32'b11110101011101011100011111010000;
   assign mem[25663:25632] = 32'b11110110000110000001100101110000;
   assign mem[25695:25664] = 32'b11111111111011100101001100011011;
   assign mem[25727:25696] = 32'b00000000110001001011110110011010;
   assign mem[25759:25728] = 32'b00000110111110110110001111010000;
   assign mem[25791:25760] = 32'b11111101011101001111000101001000;
   assign mem[25823:25792] = 32'b11111010010100000010000000001000;
   assign mem[25855:25824] = 32'b00001100011011110010000001100000;
   assign mem[25887:25856] = 32'b11111011000110001110110101110000;
   assign mem[25919:25888] = 32'b00000011101010011110010001100000;
   assign mem[25951:25920] = 32'b00000000000111001011101100000010;
   assign mem[25983:25952] = 32'b00000000111011101000000101111010;
   assign mem[26015:25984] = 32'b00000010111011100000010111011000;
   assign mem[26047:26016] = 32'b00000101001010000110001011101000;
   assign mem[26079:26048] = 32'b11111100110101101101100000100000;
   assign mem[26111:26080] = 32'b11111101010001011000110001011100;
   assign mem[26143:26112] = 32'b00000010101100110011101011100100;
   assign mem[26175:26144] = 32'b11111011000010110000000010100000;
   assign mem[26207:26176] = 32'b00000110010111011000101100101000;
   assign mem[26239:26208] = 32'b11111011000101101010011000110000;
   assign mem[26271:26240] = 32'b00000001110111011011100101111100;
   assign mem[26303:26272] = 32'b00000010110001111011101111000000;
   assign mem[26335:26304] = 32'b11111101010000010110000000100100;
   assign mem[26367:26336] = 32'b11111110010010111000101110110110;
   assign mem[26399:26368] = 32'b00000110001110011100011101001000;
   assign mem[26431:26400] = 32'b11110100000001001111001110100000;
   assign mem[26463:26432] = 32'b11111010100110111100011011000000;
   assign mem[26495:26464] = 32'b00001100101001001010001110100000;
   assign mem[26527:26496] = 32'b11111010011000011000010111010000;
   assign mem[26559:26528] = 32'b11110011011111000010111000010000;
   assign mem[26591:26560] = 32'b00000010100001111000110000000100;
   assign mem[26623:26592] = 32'b11111010001011010011011111011000;
   assign mem[26655:26624] = 32'b11111100101110100110101101010000;
   assign mem[26687:26656] = 32'b00000010010000101001101100101100;
   assign mem[26719:26688] = 32'b00000000001010001111111110001111;
   assign mem[26751:26720] = 32'b11111111110110011100001000110100;
   assign mem[26783:26752] = 32'b11110101000001011100001010100000;
   assign mem[26815:26784] = 32'b11111101001011001101101100000000;
   assign mem[26847:26816] = 32'b00000100100110010010011111111000;
   assign mem[26879:26848] = 32'b00000000101100100000011011111101;
   assign mem[26911:26880] = 32'b11111101110100010001111010100000;
   assign mem[26943:26912] = 32'b11111111001011000001011111110010;
   assign mem[26975:26944] = 32'b00000001101001111100101111000000;
   assign mem[27007:26976] = 32'b11110110100101000100010010110000;
   assign mem[27039:27008] = 32'b00000011011001100010111111111100;
   assign mem[27071:27040] = 32'b00000101010100110011101000111000;
   assign mem[27103:27072] = 32'b00001100111000101110110110010000;
   assign mem[27135:27104] = 32'b00000010100000101111100110000000;
   assign mem[27167:27136] = 32'b11111001100011011100111100001000;
   assign mem[27199:27168] = 32'b11111110011111001001100010101110;
   assign mem[27231:27200] = 32'b11111111011100101001111101000010;
   assign mem[27263:27232] = 32'b11111000111111000110101110011000;
   assign mem[27295:27264] = 32'b11111101101110100001010101100100;
   assign mem[27327:27296] = 32'b00000010111010001010101101011000;
   assign mem[27359:27328] = 32'b11110111100001000011000100000000;
   assign mem[27391:27360] = 32'b11111101111110111111110100000000;
   assign mem[27423:27392] = 32'b11110110111010001001011111100000;
   assign mem[27455:27424] = 32'b00000000001010101111010011110110;
   assign mem[27487:27456] = 32'b00000001110011100101010101111010;
   assign mem[27519:27488] = 32'b00001000100110011111001101100000;
   assign mem[27551:27520] = 32'b11110011110010100011101000100000;
   assign mem[27583:27552] = 32'b11110010101100111111100001110000;
   assign mem[27615:27584] = 32'b00000000110001001011001010000010;
   assign mem[27647:27616] = 32'b11111110001001100000101011001110;
   assign mem[27679:27648] = 32'b00000101111111011011111011011000;
   assign mem[27711:27680] = 32'b00000000101111101000001110000011;
   assign mem[27743:27712] = 32'b00000011111011011001010111110000;
   assign mem[27775:27744] = 32'b00000001010011110111011001001000;
   assign mem[27807:27776] = 32'b00000111011100110101100111010000;
   assign mem[27839:27808] = 32'b00000010010001101101001111110100;
   assign mem[27871:27840] = 32'b11110111110101110111100101000000;
   assign mem[27903:27872] = 32'b00000111000010100000101010010000;
   assign mem[27935:27904] = 32'b11111011110101110010101110100000;
   assign mem[27967:27936] = 32'b00000101111000111000010101000000;
   assign mem[27999:27968] = 32'b11111011100011101010110101010000;
   assign mem[28031:28000] = 32'b00000111110101110101011110110000;
   assign mem[28063:28032] = 32'b00000011001011011000101100010000;
   assign mem[28095:28064] = 32'b00000110010100101101110001001000;
   assign mem[28127:28096] = 32'b11111100100000111101100011000100;
   assign mem[28159:28128] = 32'b11101011011100000011010100000000;
   assign mem[28191:28160] = 32'b11101111101011101010101111000000;
   assign mem[28223:28192] = 32'b00001011110000100111000110010000;
   assign mem[28255:28224] = 32'b00000010110101000000001101000000;
   assign mem[28287:28256] = 32'b00000010001101001111111110100100;
   assign mem[28319:28288] = 32'b00001010110001000101011011110000;
   assign mem[28351:28320] = 32'b00001010010001101100010100010000;
   assign mem[28383:28352] = 32'b00000010001011001100000101100100;
   assign mem[28415:28384] = 32'b00000111001000101000111000101000;
   assign mem[28447:28416] = 32'b11110001111111111111101001100000;
   assign mem[28479:28448] = 32'b11101011011011010110010110000000;
   assign mem[28511:28480] = 32'b11110100100001010111000010000000;
   assign mem[28543:28512] = 32'b11111111010010101111011111100000;
   assign mem[28575:28544] = 32'b11110010100101000110000010110000;
   assign mem[28607:28576] = 32'b00000111011000101011101011010000;
   assign mem[28639:28608] = 32'b00000000111000010101010000000111;
   assign mem[28671:28640] = 32'b11101111101001001011001110100000;
   assign mem[28703:28672] = 32'b00010010111001100011101010000000;
   assign mem[28735:28704] = 32'b11111001100101011001100010100000;
   assign mem[28767:28736] = 32'b11111001001100111110011011001000;
   assign mem[28799:28768] = 32'b11100111100101010000100010000000;
   assign mem[28831:28800] = 32'b11110100111010100101011010110000;
   assign mem[28863:28832] = 32'b00000101011111101100011001010000;
   assign mem[28895:28864] = 32'b11101001011010101010010010000000;
   assign mem[28927:28896] = 32'b00001111100011010101000010100000;
   assign mem[28959:28928] = 32'b00000100010001101000000010011000;
   assign mem[28991:28960] = 32'b11110100100110001000110011110000;
   assign mem[29023:28992] = 32'b00001001011100111111100010100000;
   assign mem[29055:29024] = 32'b11111110100101111100101011010100;
   assign mem[29087:29056] = 32'b11111011110101010001000000111000;
   assign mem[29119:29088] = 32'b11100100101000001011011100100000;
   assign mem[29151:29120] = 32'b11111100001011110100011001000100;
   assign mem[29183:29152] = 32'b11111011101111000111100110100000;
   assign mem[29215:29184] = 32'b00000010011100111000010110110100;
   assign mem[29247:29216] = 32'b11111110111110001110011101111110;
   assign mem[29279:29248] = 32'b00000000110111000100010111000001;
   assign mem[29311:29280] = 32'b11111101110100010111011010111000;
   assign mem[29343:29312] = 32'b11111110001101001000010001111000;
   assign mem[29375:29344] = 32'b00000010100100010011100000010100;
   assign mem[29407:29376] = 32'b00000000111101000110001101000000;
   assign mem[29439:29408] = 32'b00000100000011001001101110110000;
   assign mem[29471:29440] = 32'b00000001001000001000011101100110;
   assign mem[29503:29472] = 32'b11111000100110001001100000011000;
   assign mem[29535:29504] = 32'b11111101100001011010101110010100;
   assign mem[29567:29536] = 32'b00000011000100111001111010000100;
   assign mem[29599:29568] = 32'b11110101101010010001111000100000;
   assign mem[29631:29600] = 32'b00000111000111110000101011110000;
   assign mem[29663:29632] = 32'b11111011001011011111001100001000;
   assign mem[29695:29664] = 32'b00000001000000110110001110011110;
   assign mem[29727:29696] = 32'b00000001001100001101000111100100;
   assign mem[29759:29728] = 32'b00000111111111011101011101110000;
   assign mem[29791:29760] = 32'b00000000001110011010000000101110;
   assign mem[29823:29792] = 32'b00000000011111000100100000110111;
   assign mem[29855:29824] = 32'b11111111110010100110011110000001;
   assign mem[29887:29856] = 32'b00000010010011010101011011101100;
   assign mem[29919:29888] = 32'b11111101101000000000010100100000;
   assign mem[29951:29920] = 32'b00000010100011011000111111011100;
   assign mem[29983:29952] = 32'b11110100111100011110100000100000;
   assign mem[30015:29984] = 32'b00000010110010011111010000010100;
   assign mem[30047:30016] = 32'b00000000001100110010100010101011;
   assign mem[30079:30048] = 32'b00000000111101000101111001101010;
   assign mem[30111:30080] = 32'b11111011000010011000011011101000;
   assign mem[30143:30112] = 32'b11111110100110001000000110100000;
   assign mem[30175:30144] = 32'b11110110111001011001111110010000;
   assign mem[30207:30176] = 32'b11111010111000000110101001001000;
   assign mem[30239:30208] = 32'b00001010110111000101000010100000;
   assign mem[30271:30240] = 32'b00000111101001011101001111011000;
   assign mem[30303:30272] = 32'b00001110101101110000101110000000;
   assign mem[30335:30304] = 32'b11111010100001010010111101001000;
   assign mem[30367:30336] = 32'b11111011111100000110010100001000;
   assign mem[30399:30368] = 32'b11100001101111101100101010100000;
   assign mem[30431:30400] = 32'b11101101111011101001010100100000;
   assign mem[30463:30432] = 32'b11111101101011010011001100111100;
   assign mem[30495:30464] = 32'b00000111110001011110010101010000;
   assign mem[30527:30496] = 32'b00000000100100001110111010101000;
   assign mem[30559:30528] = 32'b00000000000001001100111000101011;
   assign mem[30591:30560] = 32'b11110101111011011110010101010000;
   assign mem[30623:30592] = 32'b11111000110110100000011101110000;
   assign mem[30655:30624] = 32'b00001011100110111000000100100000;
   assign mem[30687:30656] = 32'b11111101111100010110100100010100;
   assign mem[30719:30688] = 32'b00000001100010000000010111010100;
   assign mem[30751:30720] = 32'b11110110111111100001110010010000;
   assign mem[30783:30752] = 32'b11101111000001011001000100100000;
   assign mem[30815:30784] = 32'b00000000100000000000010101010000;
   assign mem[30847:30816] = 32'b00000000001010111001100011100010;
   assign mem[30879:30848] = 32'b00000000101110101011001000011100;
   assign mem[30911:30880] = 32'b00000100100010111010111111001000;
   assign mem[30943:30912] = 32'b00000100101010101111100000000000;
   assign mem[30975:30944] = 32'b11111110101100001100100000111100;
   assign mem[31007:30976] = 32'b00000000001101110000111010000000;
   assign mem[31039:31008] = 32'b00001011111100010000100001110000;
   assign mem[31071:31040] = 32'b00000001000100100111111101001100;
   assign mem[31103:31072] = 32'b00000000100010100000000111010001;
   assign mem[31135:31104] = 32'b00000010101000111001110100000000;
   assign mem[31167:31136] = 32'b00000010001011110101011000100000;
   assign mem[31199:31168] = 32'b11111101110100001010110111000100;
   assign mem[31231:31200] = 32'b11111011101100111100101101010000;
   assign mem[31263:31232] = 32'b00000100011010001010100100000000;
   assign mem[31295:31264] = 32'b00000011011101111110000110010000;
   assign mem[31327:31296] = 32'b00001000100010111011011011010000;
   assign mem[31359:31328] = 32'b11111100110101001110100010011100;
   assign mem[31391:31360] = 32'b11111011111111110111110001111000;
   assign mem[31423:31392] = 32'b11110010010101110111111101010000;
   assign mem[31455:31424] = 32'b00000000001100000100010110001100;
   assign mem[31487:31456] = 32'b00000100111001111100111110011000;
   assign mem[31519:31488] = 32'b11101110001110111011010010100000;
   assign mem[31551:31520] = 32'b11111100001110101111011010011000;
   assign mem[31583:31552] = 32'b00000010110110000000011101100100;
   assign mem[31615:31584] = 32'b11111111010011011110010011100100;
   assign mem[31647:31616] = 32'b00000111001111111111010001010000;
   assign mem[31679:31648] = 32'b00000101010010110000011001001000;
   assign mem[31711:31680] = 32'b11111001001001001101101011010000;
   assign mem[31743:31712] = 32'b11111110001001100011010001110100;
   assign mem[31775:31744] = 32'b11111111100011001011010011000111;
   assign mem[31807:31776] = 32'b11111100111000001100011011100100;
   assign mem[31839:31808] = 32'b11111010111101010101010110000000;
   assign mem[31871:31840] = 32'b11111110101000001000101001111010;
   assign mem[31903:31872] = 32'b11111011110100100110110110011000;
   assign mem[31935:31904] = 32'b11111101001101001010000111110100;
   assign mem[31967:31936] = 32'b00000001001110011000110100000100;
   assign mem[31999:31968] = 32'b00000110001101011101000100001000;
   assign mem[32031:32000] = 32'b11111111011001111010110011001001;
   assign mem[32063:32032] = 32'b00000000100010110001110011110001;
   assign mem[32095:32064] = 32'b00000100010111010110110001010000;
   assign mem[32127:32096] = 32'b11111111100010110000110011000010;
   assign mem[32159:32128] = 32'b00000001111011111100101011110010;
   assign mem[32191:32160] = 32'b00000000000110010001110001011001;
   assign mem[32223:32192] = 32'b11110010100101100000111110000000;
   assign mem[32255:32224] = 32'b00000110001101111000000101001000;
   assign mem[32287:32256] = 32'b11111010001111001001111010000000;
   assign mem[32319:32288] = 32'b11111001101100110100101001000000;
   assign mem[32351:32320] = 32'b11111101111011000110111110101100;
   assign mem[32383:32352] = 32'b00001000001101110001100100110000;
   assign mem[32415:32384] = 32'b11111100010001101010011011110100;
   assign mem[32447:32416] = 32'b00000010011001101001010101110000;
   assign mem[32479:32448] = 32'b00001111110100010101000100110000;
   assign mem[32511:32480] = 32'b00000010100010000001000011011000;
   assign mem[32543:32512] = 32'b11111010010000101100100000010000;
   assign mem[32575:32544] = 32'b00000011011111101001011010011000;
   assign mem[32607:32576] = 32'b11111011001100010010011100110000;
   assign mem[32639:32608] = 32'b11110010010101000101010000110000;
   assign mem[32671:32640] = 32'b00000010000001111110001111100100;
   assign mem[32703:32672] = 32'b11111011000101101011100100011000;
   assign mem[32735:32704] = 32'b00000010001110011000001110111100;
   assign mem[32767:32736] = 32'b00000010101101110000100010000000;
   assign mem[32799:32768] = 32'b11111100011100110011110010110100;
   assign mem[32831:32800] = 32'b11111000111101110001110001101000;
   assign mem[32863:32832] = 32'b00001010110101011110111100100000;
   assign mem[32895:32864] = 32'b00000010011110001110010000111100;
   assign mem[32927:32896] = 32'b11111001001001011101000100010000;
   assign mem[32959:32928] = 32'b11111100010100000100111010011000;
   assign mem[32991:32960] = 32'b00000010100000100110111111000100;
   assign mem[33023:32992] = 32'b11110110001011011001001000010000;
   assign mem[33055:33024] = 32'b00000011100001100001110001111100;
   assign mem[33087:33056] = 32'b00000011101000000011011000001000;
   assign mem[33119:33088] = 32'b11111111010001010101010101111001;
   assign mem[33151:33120] = 32'b11111101111110000000111100100100;
   assign mem[33183:33152] = 32'b11111001001001110010110110101000;
   assign mem[33215:33184] = 32'b00000001000000000000100100111010;
   assign mem[33247:33216] = 32'b00000010100011011000101110111000;
   assign mem[33279:33248] = 32'b00000000110011111100100100101010;
   assign mem[33311:33280] = 32'b11110101101111111100011111110000;
   assign mem[33343:33312] = 32'b11111100000100110100110111000000;
   assign mem[33375:33344] = 32'b00001010111100000101000100110000;
   assign mem[33407:33376] = 32'b00000111010100001110000000101000;
   assign mem[33439:33408] = 32'b11110100000001010111000011100000;
   assign mem[33471:33440] = 32'b11110011000110110010001011010000;
   assign mem[33503:33472] = 32'b11111101110001011110100100001100;
   assign mem[33535:33504] = 32'b11110111110111010101100101110000;
   assign mem[33567:33536] = 32'b11111101111110001111010001101000;
   assign mem[33599:33568] = 32'b11111001111100110000010100100000;
   assign mem[33631:33600] = 32'b11110001100111110011010110000000;
   assign mem[33663:33632] = 32'b11101101001010100001110001100000;
   assign mem[33695:33664] = 32'b00000110100100111001110010111000;
   assign mem[33727:33696] = 32'b00000111000111000000110010101000;
   assign mem[33759:33728] = 32'b11110110000001101011000100010000;
   assign mem[33791:33760] = 32'b11110010111001111001000001000000;
   assign mem[33823:33792] = 32'b11111110101000100010100001111100;
   assign mem[33855:33824] = 32'b11110000101001010101011101100000;
   assign mem[33887:33856] = 32'b11111001101000011001100011100000;
   assign mem[33919:33888] = 32'b11111100011110111010100110000000;
   assign mem[33951:33920] = 32'b11110001100101000111101110010000;
   assign mem[33983:33952] = 32'b11111011101101011010111001010000;
   assign mem[34015:33984] = 32'b00001011001000010111100010010000;
   assign mem[34047:34016] = 32'b00000111100001001010111110011000;
   assign mem[34079:34048] = 32'b11111100111110000101000010111100;
   assign mem[34111:34080] = 32'b11101100111000111000100101000000;
   assign mem[34143:34112] = 32'b11111101011001000110111011111100;
   assign mem[34175:34144] = 32'b00001001101110000001011010000000;
   assign mem[34207:34176] = 32'b11111100000010000001000000110100;
   assign mem[34239:34208] = 32'b11111111000001011110110000011011;
   assign mem[34271:34240] = 32'b11111000100101011001011111100000;
   assign mem[34303:34272] = 32'b00000101010100101111001000110000;
   assign mem[34335:34304] = 32'b11111000001101110100011110101000;
   assign mem[34367:34336] = 32'b00000000100010110011101010011101;
   assign mem[34399:34368] = 32'b00001101101000101011101110110000;
   assign mem[34431:34400] = 32'b00000010001111000011001010001000;
   assign mem[34463:34432] = 32'b00001001001101001001001011100000;
   assign mem[34495:34464] = 32'b11111011100110000011100001001000;
   assign mem[34527:34496] = 32'b11110011100001111100100000100000;
   assign mem[34559:34528] = 32'b11101001011101100011101001100000;
   assign mem[34591:34560] = 32'b00000010110110100111000101100000;
   assign mem[34623:34592] = 32'b11111111011011100100100100001010;
   assign mem[34655:34624] = 32'b00000011001101111101000110011000;
   assign mem[34687:34656] = 32'b00000111000000010010111010110000;
   assign mem[34719:34688] = 32'b11110101010000110100010011100000;
   assign mem[34751:34720] = 32'b11111011101100011010111100111000;
   assign mem[34783:34752] = 32'b00000011000100001010101110001100;
   assign mem[34815:34784] = 32'b00000011010110111000110101000100;
   assign mem[34847:34816] = 32'b11110111011111100101111000100000;
   assign mem[34879:34848] = 32'b11111111111011111000100101110000;
   assign mem[34911:34880] = 32'b11111111111100010010111101001001;
   assign mem[34943:34912] = 32'b00000000101001010100011101011101;
   assign mem[34975:34944] = 32'b00000010111110111101000001101100;
   assign mem[35007:34976] = 32'b11111011011010001011101110010000;
   assign mem[35039:35008] = 32'b00000100111101111011001111011000;
   assign mem[35071:35040] = 32'b11111111100001100100110001100111;
   assign mem[35103:35072] = 32'b00000000010011011111111010010001;
   assign mem[35135:35104] = 32'b11111111011001010101000011011101;
   assign mem[35167:35136] = 32'b11111101101000111000010010000100;
   assign mem[35199:35168] = 32'b11111101001110001011101011001000;
   assign mem[35231:35200] = 32'b11111010000110001011111101010000;
   assign mem[35263:35232] = 32'b00001010110001000000110000000000;
   assign mem[35295:35264] = 32'b11111111010010010001101110010100;
   assign mem[35327:35296] = 32'b11110111100000010000010011100000;
   assign mem[35359:35328] = 32'b00000110001111111111000011100000;
   assign mem[35391:35360] = 32'b00001110010110000100000110100000;
   assign mem[35423:35392] = 32'b00000001010011001101101010011010;
   assign mem[35455:35424] = 32'b11111011011111001101001010111000;
   assign mem[35487:35456] = 32'b11111101110100000101100101110100;
   assign mem[35519:35488] = 32'b11111001000100110011101101010000;
   assign mem[35551:35520] = 32'b11111111101111011101011001011000;
   assign mem[35583:35552] = 32'b11111111110000110011010110001011;
   assign mem[35615:35584] = 32'b11111110010010100100001110010000;
   assign mem[35647:35616] = 32'b00000010010000010000011001010100;
   assign mem[35679:35648] = 32'b00000001111101001111001000010010;
   assign mem[35711:35680] = 32'b11111100101100100101111101100100;
   assign mem[35743:35712] = 32'b00000000010001111100111100011001;
   assign mem[35775:35744] = 32'b00000001011011100100110010001110;
   assign mem[35807:35776] = 32'b00000000111100011011001001001001;
   assign mem[35839:35808] = 32'b00000001010011110111111011011010;
   assign mem[35871:35840] = 32'b00000110101110001001010111000000;
   assign mem[35903:35872] = 32'b11101110001010100001111100100000;
   assign mem[35935:35904] = 32'b00000111100011110110101011011000;
   assign mem[35967:35936] = 32'b11111010001110100111110000010000;
   assign mem[35999:35968] = 32'b11110110100100111101001100110000;
   assign mem[36031:36000] = 32'b11111100011001111110011110110100;
   assign mem[36063:36032] = 32'b00001000100011011011000010110000;
   assign mem[36095:36064] = 32'b11111100101010011001000010101000;
   assign mem[36127:36096] = 32'b11111111000010001100111110001001;
   assign mem[36159:36128] = 32'b00000000000101011010010101100000;
   assign mem[36191:36160] = 32'b00000001001000010111101010000110;
   assign mem[36223:36192] = 32'b11111101100011001100001110111100;
   assign mem[36255:36224] = 32'b00000100001010010000110111011000;
   assign mem[36287:36256] = 32'b11111011111110101000000101001000;
   assign mem[36319:36288] = 32'b00000000111110010110001110010010;
   assign mem[36351:36320] = 32'b11111111110111111011101110011000;
   assign mem[36383:36352] = 32'b11111111011100101010001100010101;
   assign mem[36415:36384] = 32'b11111101110000110110010011010000;
   assign mem[36447:36416] = 32'b00000101000000000110000001000000;
   assign mem[36479:36448] = 32'b11111110001100011010001110010010;
   assign mem[36511:36480] = 32'b11111101111111110011011110000000;
   assign mem[36543:36512] = 32'b11111111000101010010011111110111;
   assign mem[36575:36544] = 32'b00000000010110111000100001110100;
   assign mem[36607:36576] = 32'b00000010010111000010100000101000;
   assign mem[36639:36608] = 32'b11110111001110000001010101010000;
   assign mem[36671:36640] = 32'b11111000011001011101100011110000;
   assign mem[36703:36672] = 32'b00000101110001111011001111011000;
   assign mem[36735:36704] = 32'b11111011010001111000011101010000;
   assign mem[36767:36736] = 32'b00001010100111011111000000110000;
   assign mem[36799:36768] = 32'b00001011010110111001110001010000;
   assign mem[36831:36800] = 32'b11110111001010001111110001100000;
   assign mem[36863:36832] = 32'b00000011010001001000010000111000;
   assign mem[36895:36864] = 32'b11111101110010000011000010100100;
   assign mem[36927:36896] = 32'b00000010010111011000111111011000;
   assign mem[36959:36928] = 32'b00000110000111100101011011000000;
   assign mem[36991:36960] = 32'b11111110111100010110011110000010;
   assign mem[37023:36992] = 32'b11111010110011001111111010000000;
   assign mem[37055:37024] = 32'b00000000001000110011100111101111;
   assign mem[37087:37056] = 32'b00000110110010010101001101000000;
   assign mem[37119:37088] = 32'b11111110001100000100011101110000;
   assign mem[37151:37120] = 32'b11110010111111110000100101100000;
   assign mem[37183:37152] = 32'b11111111000110001101100001100100;
   assign mem[37215:37184] = 32'b00000000111100110000110001101110;
   assign mem[37247:37216] = 32'b00000011111001010010000100111000;
   assign mem[37279:37248] = 32'b11111010011111100011001011000000;
   assign mem[37311:37280] = 32'b11111110001101110110111010000010;
   assign mem[37343:37312] = 32'b11111101011101111001100011111100;
   assign mem[37375:37344] = 32'b00000111100000100111101000101000;
   assign mem[37407:37376] = 32'b00000011110010010000010010110100;
   assign mem[37439:37408] = 32'b00000000010111010111111000110101;
   assign mem[37471:37440] = 32'b00000000111011100111110000000100;
   assign mem[37503:37472] = 32'b11110101101011111101100100000000;
   assign mem[37535:37504] = 32'b00000011011000010111001001000100;
   assign mem[37567:37536] = 32'b00000000111100111110111011100000;
   assign mem[37599:37568] = 32'b11110100000001111111010111110000;
   assign mem[37631:37600] = 32'b00000100000110010000100011000000;
   assign mem[37663:37632] = 32'b00000010011011011100010111001100;
   assign mem[37695:37664] = 32'b00000100100011000010100111110000;
   assign mem[37727:37696] = 32'b00000000001010010000001101101001;
   assign mem[37759:37728] = 32'b00000001100100001110010001100110;
   assign mem[37791:37760] = 32'b11110101010001111111100111000000;
   assign mem[37823:37792] = 32'b11110100111010001110101010100000;
   assign mem[37855:37824] = 32'b00001000011110010110111100010000;
   assign mem[37887:37856] = 32'b00000011011001111000100010000100;
   assign mem[37919:37888] = 32'b11110101000111010111001100100000;
   assign mem[37951:37920] = 32'b11111110111110010111111100011100;
   assign mem[37983:37952] = 32'b00000011011100001100111101100100;
   assign mem[38015:37984] = 32'b00000010001110011101111100011100;
   assign mem[38047:38016] = 32'b11111110101111011011010001011100;
   assign mem[38079:38048] = 32'b00000101111010001100111010001000;
   assign mem[38111:38080] = 32'b11111011011011110110001100110000;
   assign mem[38143:38112] = 32'b00000010111101111111101010011100;
   assign mem[38175:38144] = 32'b11111011000010101011101101111000;
   assign mem[38207:38176] = 32'b11111101011001001001111001101000;
   assign mem[38239:38208] = 32'b00000011010101101101111101011000;
   assign mem[38271:38240] = 32'b00000111011000010111100110110000;
   assign mem[38303:38272] = 32'b00001010101000101010010110100000;
   assign mem[38335:38304] = 32'b11111101010001101111100011100000;
   assign mem[38367:38336] = 32'b11111100010101010111100100110000;
   assign mem[38399:38368] = 32'b11110101011000101101111000010000;
   assign mem[38431:38400] = 32'b11110111111111000010101100010000;
   assign mem[38463:38432] = 32'b11111111000100100110011100000100;
   assign mem[38495:38464] = 32'b11111110001110010001111111101000;
   assign mem[38527:38496] = 32'b11111111000111011010110011100000;
   assign mem[38559:38528] = 32'b00000010100010110111110000011000;
   assign mem[38591:38560] = 32'b11111001011110100110111010110000;
   assign mem[38623:38592] = 32'b11111111100101011101110111010111;
   assign mem[38655:38624] = 32'b11111111111100010110110000001011;
   assign mem[38687:38656] = 32'b00001000011001010111111101110000;
   assign mem[38719:38688] = 32'b11110100111100001101101010110000;
   assign mem[38751:38720] = 32'b11111001111111110111011000001000;
   assign mem[38783:38752] = 32'b00000010100011110010000000010000;
   assign mem[38815:38784] = 32'b00000101111011001000111000101000;
   assign mem[38847:38816] = 32'b00001001011100011011100111100000;
   assign mem[38879:38848] = 32'b11111011110111100101011001111000;
   assign mem[38911:38880] = 32'b11110110111010000110000110000000;
   assign mem[38943:38912] = 32'b11111100011000101101111110100100;
   assign mem[38975:38944] = 32'b00000101000001000110111001100000;
   assign mem[39007:38976] = 32'b11111011000101011000001100101000;
   assign mem[39039:39008] = 32'b11101001001101001001110101000000;
   assign mem[39071:39040] = 32'b11111011110111110101110110010000;
   assign mem[39103:39072] = 32'b11111100110100001001100011100100;
   assign mem[39135:39104] = 32'b00000000111010000111110101110110;
   assign mem[39167:39136] = 32'b00000001011000000011101111111010;
   assign mem[39199:39168] = 32'b11111111111001000011111110010010;
   assign mem[39231:39200] = 32'b11111011100001011010011000110000;
   assign mem[39263:39232] = 32'b11111100001011000110011111111000;
   assign mem[39295:39264] = 32'b00000010111100001001011110111000;
   assign mem[39327:39296] = 32'b00000011010111011111111001111100;
   assign mem[39359:39328] = 32'b00000001000010011100100110000100;
   assign mem[39391:39360] = 32'b11111011010101111000000111000000;
   assign mem[39423:39392] = 32'b00000001010110101101000101101100;
   assign mem[39455:39424] = 32'b11111111001011110011101100011001;
   assign mem[39487:39456] = 32'b11111110111001001000101000101110;
   assign mem[39519:39488] = 32'b11111110100100110011001000011100;
   assign mem[39551:39520] = 32'b00000011100110001110101010110100;
   assign mem[39583:39552] = 32'b00000000101111101100011000110101;
   assign mem[39615:39584] = 32'b00000011010110101000001111111000;
   assign mem[39647:39616] = 32'b00000000010010011101100100001100;
   assign mem[39679:39648] = 32'b11111111101111100010001011010010;
   assign mem[39711:39680] = 32'b00000000010110010100000001101000;
   assign mem[39743:39712] = 32'b11111101011101010111111011101000;
   assign mem[39775:39744] = 32'b11111111011000010100111011100000;
   assign mem[39807:39776] = 32'b00000000011001100110000110111010;
   assign mem[39839:39808] = 32'b00000000100000000111110001011101;
   assign mem[39871:39840] = 32'b11111111100111101101100111101011;
   assign mem[39903:39872] = 32'b11110111111001000000011001110000;
   assign mem[39935:39904] = 32'b11111110110000101101011010100010;
   assign mem[39967:39936] = 32'b00000000100000101010000101100010;
   assign mem[39999:39968] = 32'b11111101101000101100001000011100;
   assign mem[40031:40000] = 32'b11111101011101011100111101001000;
   assign mem[40063:40032] = 32'b11111011111000100001001001111000;
   assign mem[40095:40064] = 32'b00000001101110100011011111010110;
   assign mem[40127:40096] = 32'b11111111001110010000000000110000;
   assign mem[40159:40128] = 32'b11111110101101010100101110101000;
   assign mem[40191:40160] = 32'b11111100110110110011111101011000;
   assign mem[40223:40192] = 32'b00000001001101000100110100101100;
   assign mem[40255:40224] = 32'b11111100000010011010000000100100;
   assign mem[40287:40256] = 32'b00000111011110001011111001010000;
   assign mem[40319:40288] = 32'b11111111000111010100100001001011;
   assign mem[40351:40320] = 32'b11111111000000101101100101111001;
   assign mem[40383:40352] = 32'b00000100110000000101100011110000;
   assign mem[40415:40384] = 32'b00000001001111110100011100011100;
   assign mem[40447:40416] = 32'b11111011100000000010011101011000;
   assign mem[40479:40448] = 32'b00000011100011110000010011110000;
   assign mem[40511:40480] = 32'b00000000101010011001111010111011;
   assign mem[40543:40512] = 32'b00000000001011000110100010111001;
   assign mem[40575:40544] = 32'b00000000001000111110011100000010;
   assign mem[40607:40576] = 32'b00000100011001100101101101111000;
   assign mem[40639:40608] = 32'b11111101011010010000011010000000;
   assign mem[40671:40640] = 32'b11111111100010001001110100011100;
   assign mem[40703:40672] = 32'b00000110010101101111111000110000;
   assign mem[40735:40704] = 32'b11111100000101111000000110110000;
   assign mem[40767:40736] = 32'b11110110011011000010111100010000;
   assign mem[40799:40768] = 32'b00000010101010100011100100001100;
   assign mem[40831:40800] = 32'b00000011110000000111011111111100;
   assign mem[40863:40832] = 32'b00000110001000001101111010011000;
   assign mem[40895:40864] = 32'b00000011010011011100000101010000;
   assign mem[40927:40896] = 32'b11111100110001101110100100101100;
   assign mem[40959:40928] = 32'b11111011100111000011000011010000;
   assign mem[40991:40960] = 32'b11111001011101100101010110101000;
   assign mem[41023:40992] = 32'b11101111110001010000011001000000;
   assign mem[41055:41024] = 32'b00000010000000100010110001000100;
   assign mem[41087:41056] = 32'b00000101010100000010011111010000;
   assign mem[41119:41088] = 32'b11111011001011110010111100101000;
   assign mem[41151:41120] = 32'b00000011010001111101100100101000;
   assign mem[41183:41152] = 32'b11110011000101100101100101000000;
   assign mem[41215:41184] = 32'b00000011101011000110011101110000;
   assign mem[41247:41216] = 32'b11111110011010001100101000011110;
   assign mem[41279:41248] = 32'b00000000101100010110100100001111;
   assign mem[41311:41280] = 32'b11111010110001000100010010100000;
   assign mem[41343:41312] = 32'b00000010011110101110010100100100;
   assign mem[41375:41344] = 32'b00000011110010011001100001011000;
   assign mem[41407:41376] = 32'b00000010111010100100111011101100;
   assign mem[41439:41408] = 32'b00001001111011110001011100100000;
   assign mem[41471:41440] = 32'b11110010101011110110110010110000;
   assign mem[41503:41472] = 32'b00000000010110000100010100001100;
   assign mem[41535:41504] = 32'b00000101101000100011011000111000;
   assign mem[41567:41536] = 32'b11110111110100110101000111110000;
   assign mem[41599:41568] = 32'b11110111011101101010011000110000;
   assign mem[41631:41600] = 32'b00000100111000001100010100111000;
   assign mem[41663:41632] = 32'b11110111110011011110011011110000;
   assign mem[41695:41664] = 32'b00000110111000011101100000011000;
   assign mem[41727:41696] = 32'b00000000010101000001001100101011;
   assign mem[41759:41728] = 32'b11110101000111100001010100110000;
   assign mem[41791:41760] = 32'b11111000001110110011010011100000;
   assign mem[41823:41792] = 32'b11111111001010011000001110001110;
   assign mem[41855:41824] = 32'b11111111011110110101101100101100;
   assign mem[41887:41856] = 32'b00000011110110101101011111011100;
   assign mem[41919:41888] = 32'b00000101101110001011110001101000;
   assign mem[41951:41920] = 32'b11111000001001100101010001101000;
   assign mem[41983:41952] = 32'b11111011110111000010001011111000;
   assign mem[42015:41984] = 32'b00000010000011000100010110100100;
   assign mem[42047:42016] = 32'b00001011111101100111000010010000;
   assign mem[42079:42048] = 32'b11110111111110100000011101010000;
   assign mem[42111:42080] = 32'b11110011000101111011111100100000;
   assign mem[42143:42112] = 32'b11111010110010010110101100110000;
   assign mem[42175:42144] = 32'b00000010011000011101101100001000;
   assign mem[42207:42176] = 32'b11111101011101101000010011010100;
   assign mem[42239:42208] = 32'b00000101110110101101101100000000;
   assign mem[42271:42240] = 32'b00000101001011100100100010111000;
   assign mem[42303:42272] = 32'b11111000001001101110000000111000;
   assign mem[42335:42304] = 32'b00000011101010000110111110001100;
   assign mem[42367:42336] = 32'b00000010000000000101001001110000;
   assign mem[42399:42368] = 32'b11101110001010010010010101000000;
   assign mem[42431:42400] = 32'b11111001000100000011010001001000;
   assign mem[42463:42432] = 32'b00000001100001011101011110010010;
   assign mem[42495:42464] = 32'b11110011111111001100110111010000;
   assign mem[42527:42496] = 32'b11111100010011101110011101100000;
   assign mem[42559:42528] = 32'b00000100100111100000011001001000;
   assign mem[42591:42560] = 32'b00000111010011000110010111000000;
   assign mem[42623:42592] = 32'b00000111111000000010100101110000;
   assign mem[42655:42624] = 32'b11111011111101100001110111010000;
   assign mem[42687:42656] = 32'b11111100100101111100000010111100;
   assign mem[42719:42688] = 32'b11111001010001111010111000110000;
   assign mem[42751:42720] = 32'b11111110001001001111010011000110;
   assign mem[42783:42752] = 32'b11111110110100111111000101111110;
   assign mem[42815:42784] = 32'b00000001110010010110001110111000;
   assign mem[42847:42816] = 32'b00000011111011010000101000101100;
   assign mem[42879:42848] = 32'b00000011111001010111101111010100;
   assign mem[42911:42880] = 32'b11101111100101101100010011100000;
   assign mem[42943:42912] = 32'b00001101011001010001110110000000;
   assign mem[42975:42944] = 32'b11110110001101001010001010110000;
   assign mem[43007:42976] = 32'b11110000010000101100100111010000;
   assign mem[43039:43008] = 32'b00001010011111001100001000000000;
   assign mem[43071:43040] = 32'b11111101100000110101011101010000;
   assign mem[43103:43072] = 32'b00011010000110100011110000000000;
   assign mem[43135:43104] = 32'b11101101100010111001010101100000;
   assign mem[43167:43136] = 32'b11111100011110111110001100001000;
   assign mem[43199:43168] = 32'b11101001100100011011110000100000;
   assign mem[43231:43200] = 32'b11111111001000101010110000111000;
   assign mem[43263:43232] = 32'b00001010010010010100110110110000;
   assign mem[43295:43264] = 32'b11111011101010101011010101101000;
   assign mem[43327:43296] = 32'b11111010100100101011011101100000;
   assign mem[43359:43328] = 32'b00000000000101011011110100001011;
   assign mem[43391:43360] = 32'b00000100100111111000011011011000;
   assign mem[43423:43392] = 32'b00000011000000011011110000011000;
   assign mem[43455:43424] = 32'b11101000001110001111011101000000;
   assign mem[43487:43456] = 32'b00000111010011111110010000000000;
   assign mem[43519:43488] = 32'b11111010011110111100010111010000;
   assign mem[43551:43520] = 32'b00000100011011011110000001011000;
   assign mem[43583:43552] = 32'b00000000111001001011100101111000;
   assign mem[43615:43584] = 32'b11111111101100110000111001010010;
   assign mem[43647:43616] = 32'b00000001010010010101011101001100;
   assign mem[43679:43648] = 32'b00000001011010010101100001001000;
   assign mem[43711:43680] = 32'b11111101110111111101100011000100;
   assign mem[43743:43712] = 32'b11111000011100100111101000011000;
   assign mem[43775:43744] = 32'b00000011101100010110010000001100;
   assign mem[43807:43776] = 32'b00000000111000100000010010011100;
   assign mem[43839:43808] = 32'b00000010111110100001011101001100;
   assign mem[43871:43840] = 32'b11111111001101101001011101000010;
   assign mem[43903:43872] = 32'b00000011011010000111001001010100;
   assign mem[43935:43904] = 32'b11111011010101011100011100110000;
   assign mem[43967:43936] = 32'b11111001110010110110110000010000;
   assign mem[43999:43968] = 32'b00001000110000001100100000010000;
   assign mem[44031:44000] = 32'b00000010101100010110011011000000;
   assign mem[44063:44032] = 32'b00000110000100100111000001011000;
   assign mem[44095:44064] = 32'b11110010000011011011011101100000;
   assign mem[44127:44096] = 32'b11111010000110101101001111111000;
   assign mem[44159:44128] = 32'b11111000010011111100010110110000;
   assign mem[44191:44160] = 32'b11111001011111110010110101111000;
   assign mem[44223:44192] = 32'b11110110100010110011001111010000;
   assign mem[44255:44224] = 32'b11111111010100111110010000101100;
   assign mem[44287:44256] = 32'b00000001011100111111101010001100;
   assign mem[44319:44288] = 32'b11110111101000011101111100010000;
   assign mem[44351:44320] = 32'b11111110111011010001011110010110;
   assign mem[44383:44352] = 32'b11111101010011011100010100111100;
   assign mem[44415:44384] = 32'b00000000101111001110101101001000;
   assign mem[44447:44416] = 32'b00000010011111101100100010010000;
   assign mem[44479:44448] = 32'b00000011010110111101111111110000;
   assign mem[44511:44480] = 32'b11111001101111101100000011011000;
   assign mem[44543:44512] = 32'b00000110110001001011011001001000;
   assign mem[44575:44544] = 32'b00000011101010001001000110011000;
   assign mem[44607:44576] = 32'b00000100010001100010101110010000;
   assign mem[44639:44608] = 32'b00000001110110001000100011110000;
   assign mem[44671:44640] = 32'b11110011101101010101000101010000;
   assign mem[44703:44672] = 32'b11111111000110101010001001110000;
   assign mem[44735:44704] = 32'b11111110101101000011000111011110;
   assign mem[44767:44736] = 32'b00000100000100011000000110011000;
   assign mem[44799:44768] = 32'b11110011100100010011111111010000;
   assign mem[44831:44800] = 32'b11111110000100110110011101110100;
   assign mem[44863:44832] = 32'b11111011111010011000101000111000;
   assign mem[44895:44864] = 32'b00000000111000111011011110111011;
   assign mem[44927:44896] = 32'b00000010011011011001000100001100;
   assign mem[44959:44928] = 32'b11110010110000101001100011000000;
   assign mem[44991:44960] = 32'b00000000111110011011001010011100;
   assign mem[45023:44992] = 32'b11111000000101001100011110111000;
   assign mem[45055:45024] = 32'b00000001001010010000011100001100;
   assign mem[45087:45056] = 32'b00000000101110010110011010100000;
   assign mem[45119:45088] = 32'b00000010010110010011001010011000;
   assign mem[45151:45120] = 32'b11111111000010011111010110110010;
   assign mem[45183:45152] = 32'b11111010110100110110010100011000;
   assign mem[45215:45184] = 32'b11111111100011100101100101011011;
   assign mem[45247:45216] = 32'b00000000001011110010100000000011;
   assign mem[45279:45248] = 32'b11111001011100110100110100010000;
   assign mem[45311:45280] = 32'b11111100110110100111000000011000;
   assign mem[45343:45312] = 32'b11110101101101101110111000000000;
   assign mem[45375:45344] = 32'b00000011110000010100000100001000;
   assign mem[45407:45376] = 32'b00000000000111000000010101011100;
   assign mem[45439:45408] = 32'b00000011101110011101011111010100;
   assign mem[45471:45440] = 32'b00000001001101011111010101010110;
   assign mem[45503:45472] = 32'b11110111011011001010001101110000;
   assign mem[45535:45504] = 32'b00000000100010000100101111010111;
   assign mem[45567:45536] = 32'b00000100100000011011111110010000;
   assign mem[45599:45568] = 32'b11110010111111100001001100010000;
   assign mem[45631:45600] = 32'b00000100100101100011011100011000;
   assign mem[45663:45632] = 32'b11111001011100110001000001111000;
   assign mem[45695:45664] = 32'b00000110000001110110110011000000;
   assign mem[45727:45696] = 32'b11111100100110101110001101000000;
   assign mem[45759:45728] = 32'b11111010011101000101111001000000;
   assign mem[45791:45760] = 32'b00000001000000000001010100111110;
   assign mem[45823:45792] = 32'b00000000110111010001100001111100;
   assign mem[45855:45824] = 32'b11111110000011001111101011001110;
   assign mem[45887:45856] = 32'b11111011010101110100010100100000;
   assign mem[45919:45888] = 32'b00000000011100100011111010010101;
   assign mem[45951:45920] = 32'b00000011110011101110000110111100;
   assign mem[45983:45952] = 32'b00000100010101010110011010011000;
   assign mem[46015:45984] = 32'b11110101111100101000000100110000;
   assign mem[46047:46016] = 32'b11111111110011011000111101100011;
   assign mem[46079:46048] = 32'b11111110110001101101000101111100;
   assign mem[46111:46080] = 32'b11111101110011010111011110100100;
   assign mem[46143:46112] = 32'b00000000100101110000000110001101;
   assign mem[46175:46144] = 32'b11111110111000010111000011001000;
   assign mem[46207:46176] = 32'b11111111001010000001101100100101;
   assign mem[46239:46208] = 32'b11110100110000111101110000100000;
   assign mem[46271:46240] = 32'b00000110001010011001000000100000;
   assign mem[46303:46272] = 32'b11111001100001100010001001100000;
   assign mem[46335:46304] = 32'b00000011010100000011110010111000;
   assign mem[46367:46336] = 32'b11111110110001000001100010100010;
   assign mem[46399:46368] = 32'b11111110001010101001100011111010;
   assign mem[46431:46400] = 32'b11111001000100111011011110111000;
   assign mem[46463:46432] = 32'b11111101100100100011011011110100;
   assign mem[46495:46464] = 32'b00000011010000111111000000111000;
   assign mem[46527:46496] = 32'b00000000011011000011100001001101;
   assign mem[46559:46528] = 32'b11110110000101101111111100100000;
   assign mem[46591:46560] = 32'b11111110000101110011110010110010;
   assign mem[46623:46592] = 32'b11110111100010001100101010010000;
   assign mem[46655:46624] = 32'b11111110100111000101100000000010;
   assign mem[46687:46656] = 32'b00000010111011011000011001000000;
   assign mem[46719:46688] = 32'b00000010111100110111100101010100;
   assign mem[46751:46720] = 32'b11111110110010101011101100101000;
   assign mem[46783:46752] = 32'b11111101010110100001101111001100;
   assign mem[46815:46784] = 32'b00000100010001100010101011101000;
   assign mem[46847:46816] = 32'b00000100010000000010000111101000;
   assign mem[46879:46848] = 32'b00000111000001000111100001110000;
   assign mem[46911:46880] = 32'b00000000100110011011011110010110;
   assign mem[46943:46912] = 32'b11110101001001101010101100110000;
   assign mem[46975:46944] = 32'b00000110001000001100111110110000;
   assign mem[47007:46976] = 32'b11111000000111101101101000100000;
   assign mem[47039:47008] = 32'b11111110000100111101101010011110;
   assign mem[47071:47040] = 32'b11111101100110110010111011000000;
   assign mem[47103:47072] = 32'b00000001100000110100001010100100;
   assign mem[47135:47104] = 32'b00000100101100110111000110110000;
   assign mem[47167:47136] = 32'b00000001101111100010010000011010;
   assign mem[47199:47168] = 32'b11111010100011101100010111111000;
   assign mem[47231:47200] = 32'b00000001001011110100111011111110;
   assign mem[47263:47232] = 32'b11111010111110111110011001101000;
   assign mem[47295:47264] = 32'b11111110011111001001001010101010;
   assign mem[47327:47296] = 32'b00000010011111001011000011101000;
   assign mem[47359:47328] = 32'b00001000111010100101011010100000;
   assign mem[47391:47360] = 32'b11111010011011001011001011001000;
   assign mem[47423:47392] = 32'b00000101010001101011100000010000;
   assign mem[47455:47424] = 32'b11111010001100100101111101011000;
   assign mem[47487:47456] = 32'b11110110100101011101111110100000;
   assign mem[47519:47488] = 32'b00000100101101100111001100001000;
   assign mem[47551:47520] = 32'b00001000011100111111110010100000;
   assign mem[47583:47552] = 32'b00000100100011110110000111001000;
   assign mem[47615:47584] = 32'b11111000111001001001000101111000;
   assign mem[47647:47616] = 32'b00000001011100001011110011101100;
   assign mem[47679:47648] = 32'b11110101000111101001001101100000;
   assign mem[47711:47680] = 32'b11111011100000001100111110010000;
   assign mem[47743:47712] = 32'b11111001111011101100111001000000;
   assign mem[47775:47744] = 32'b11111111001001001111100110010101;
   assign mem[47807:47776] = 32'b00000001101001111110010010010100;
   assign mem[47839:47808] = 32'b11110111111110000111110111100000;
   assign mem[47871:47840] = 32'b11111110100001100000111101000000;
   assign mem[47903:47872] = 32'b11111111111000000100101100100001;
   assign mem[47935:47904] = 32'b00000000011100000000001110000110;
   assign mem[47967:47936] = 32'b00000001111000010100110011110010;
   assign mem[47999:47968] = 32'b00000110101000101011000001001000;
   assign mem[48031:48000] = 32'b00000001000011001001010110100010;
   assign mem[48063:48032] = 32'b00000100001111111001011101001000;
   assign mem[48095:48064] = 32'b00000001010111111111101001001010;
   assign mem[48127:48096] = 32'b11110110000011101101110011010000;
   assign mem[48159:48128] = 32'b00000100100000111111100011111000;
   assign mem[48191:48160] = 32'b11111111011110001000001010000010;
   assign mem[48223:48192] = 32'b11111110010011010001010001101100;
   assign mem[48255:48224] = 32'b11110100110110100001000010000000;
   assign mem[48287:48256] = 32'b11111111111100101001110111110101;
   assign mem[48319:48288] = 32'b00000001100101100000011011001110;
   assign mem[48351:48320] = 32'b11111111110001100101011000100001;
   assign mem[48383:48352] = 32'b00000101010010010100001000111000;
   assign mem[48415:48384] = 32'b00000101110111110110000010010000;
   assign mem[48447:48416] = 32'b00000000001000101001110000101001;
   assign mem[48479:48448] = 32'b00000100001101010001101100001000;
   assign mem[48511:48480] = 32'b11111111100001101001001101000011;
   assign mem[48543:48512] = 32'b11111100000101111110100101100100;
   assign mem[48575:48544] = 32'b00000101101010001011111000000000;
   assign mem[48607:48576] = 32'b11111000110101110101101001010000;
   assign mem[48639:48608] = 32'b11110010010111001111110001110000;
   assign mem[48671:48640] = 32'b11111101101101101111011001001000;
   assign mem[48703:48672] = 32'b00001100101010111100010100000000;
   assign mem[48735:48704] = 32'b00000010011000101100001011000000;
   assign mem[48767:48736] = 32'b11111110110000001110001010001110;
   assign mem[48799:48768] = 32'b00000101110111010000000110111000;
   assign mem[48831:48800] = 32'b00000000101110001010101100011010;
   assign mem[48863:48832] = 32'b11111110001010000011111101010010;
   assign mem[48895:48864] = 32'b11111110111001000101101100010110;
   assign mem[48927:48896] = 32'b11111101010100001010011110001100;
   assign mem[48959:48928] = 32'b11110010111000000110111100010000;
   assign mem[48991:48960] = 32'b11110110111001111111010000010000;
   assign mem[49023:48992] = 32'b00001100101001000110111000100000;
   assign mem[49055:49024] = 32'b00000001011101101011101011100110;
   assign mem[49087:49056] = 32'b00001010011010100110000111010000;
   assign mem[49119:49088] = 32'b00001001111111111100111010010000;
   assign mem[49151:49120] = 32'b11101001000000110101101100000000;
   assign mem[49183:49152] = 32'b00001110110110001011001101110000;
   assign mem[49215:49184] = 32'b11101001101111111000110110100000;
   assign mem[49247:49216] = 32'b11111100011100000111010110100100;
   assign mem[49279:49248] = 32'b11100101100000101110100111100000;
   assign mem[49311:49280] = 32'b11110100111111000011110100110000;
   assign mem[49343:49312] = 32'b00001011111000110000010100100000;
   assign mem[49375:49344] = 32'b11111110011111001111010010111010;
   assign mem[49407:49376] = 32'b11111111111101001000101011010100;
   assign mem[49439:49408] = 32'b00001000100101100010001101000000;
   assign mem[49471:49440] = 32'b11111100111010001111100101110100;
   assign mem[49503:49472] = 32'b00001001000011110001100000010000;
   assign mem[49535:49504] = 32'b00000110000000010101101010101000;
   assign mem[49567:49536] = 32'b11110100001111101100010011110000;
   assign mem[49599:49568] = 32'b11100110100110001110000100000000;
   assign mem[49631:49600] = 32'b00000011011110100111011101000000;
   assign mem[49663:49632] = 32'b00000100110101011110011001010000;
   assign mem[49695:49664] = 32'b11111110101101000100001100101000;
   assign mem[49727:49696] = 32'b11111100001110111001001111011000;
   assign mem[49759:49728] = 32'b00000000010100100110101110011010;
   assign mem[49791:49760] = 32'b00000000101000001111100101111100;
   assign mem[49823:49792] = 32'b00000100001001000101110000110000;
   assign mem[49855:49824] = 32'b11111110000010011111001000000110;
   assign mem[49887:49856] = 32'b00000001110110001111100000001010;
   assign mem[49919:49888] = 32'b00000000011001011101100011110011;
   assign mem[49951:49920] = 32'b11111011011000011010100011100000;
   assign mem[49983:49952] = 32'b11111101101001010101000111000100;
   assign mem[50015:49984] = 32'b11111110011011100011010011110110;
   assign mem[50047:50016] = 32'b00000001001011101111110011011000;
   assign mem[50079:50048] = 32'b11110011000001010001101100010000;
   assign mem[50111:50080] = 32'b00000100101011011110011011111000;
   assign mem[50143:50112] = 32'b11110111111101101001000010010000;
   assign mem[50175:50144] = 32'b00000101010000011111000111101000;
   assign mem[50207:50176] = 32'b11111111100111010011001110000010;
   assign mem[50239:50208] = 32'b00000010110110111001001011001100;
   assign mem[50271:50240] = 32'b11111111011110010101011101010110;
   assign mem[50303:50272] = 32'b11111101000001110011001100100000;
   assign mem[50335:50304] = 32'b00000010110101111110010100011100;
   assign mem[50367:50336] = 32'b00000100100101100110001001001000;
   assign mem[50399:50368] = 32'b11111100100001000101001000111000;
   assign mem[50431:50400] = 32'b00000001110000101001111010000110;
   assign mem[50463:50432] = 32'b11111001111101111010111000011000;
   assign mem[50495:50464] = 32'b00000010111010011100111101011100;
   assign mem[50527:50496] = 32'b00000011010000010100111001101100;
   assign mem[50559:50528] = 32'b00000011010111110000010010001100;
   assign mem[50591:50560] = 32'b11110111010001100011011101010000;
   assign mem[50623:50592] = 32'b00010000010000001000100101000000;
   assign mem[50655:50624] = 32'b11110111110000110111010001000000;
   assign mem[50687:50656] = 32'b11110111100101001101011010000000;
   assign mem[50719:50688] = 32'b00010001001010101101010001000000;
   assign mem[50751:50720] = 32'b00000111011101100110110100001000;
   assign mem[50783:50752] = 32'b00001101100100110100011110110000;
   assign mem[50815:50784] = 32'b00000111010100010100100111010000;
   assign mem[50847:50816] = 32'b11110100010110011010110010000000;
   assign mem[50879:50848] = 32'b11101000000010111111011110100000;
   assign mem[50911:50880] = 32'b11111110001111110110101101110000;
   assign mem[50943:50912] = 32'b11111101100011000000111100000100;
   assign mem[50975:50944] = 32'b00000001101000101011010100111010;
   assign mem[51007:50976] = 32'b00000000000101011111001001001010;
   assign mem[51039:51008] = 32'b11101001101000000000101100000000;
   assign mem[51071:51040] = 32'b00000010111011011110000100001100;
   assign mem[51103:51072] = 32'b11111000000111100111011011010000;
   assign mem[51135:51104] = 32'b00001001000000001100001011000000;
   assign mem[51167:51136] = 32'b00000010000110000000011100110100;
   assign mem[51199:51168] = 32'b00000000111110001000111001010001;
   assign mem[51231:51200] = 32'b00000010011110110010101001111000;
   assign mem[51263:51232] = 32'b00001001011110001111011111110000;
   assign mem[51295:51264] = 32'b00000010100010110010000101010000;
   assign mem[51327:51296] = 32'b00000001000011111101111100001000;
   assign mem[51359:51328] = 32'b11111001111110001001010110001000;
   assign mem[51391:51360] = 32'b00000011101110101101101000001000;
   assign mem[51423:51392] = 32'b11111111111011100000110111011100;
   assign mem[51455:51424] = 32'b11111001100001010110001110001000;
   assign mem[51487:51456] = 32'b11111110101100010000101001101000;
   assign mem[51519:51488] = 32'b11110111101111001100010111000000;
   assign mem[51551:51520] = 32'b11111101110010001000110111010100;
   assign mem[51583:51552] = 32'b00000011000100100101100000000100;
   assign mem[51615:51584] = 32'b00000001000111110001110000110000;
   assign mem[51647:51616] = 32'b11111101000111111111000000101000;
   assign mem[51679:51648] = 32'b00001010010011101000010111000000;
   assign mem[51711:51680] = 32'b00000000100001001101000011111000;
   assign mem[51743:51712] = 32'b00000010101101001101101001000000;
   assign mem[51775:51744] = 32'b11110001001101010100110011100000;
   assign mem[51807:51776] = 32'b11111111011100000101100100010001;
   assign mem[51839:51808] = 32'b11111011100011110001000101000000;
   assign mem[51871:51840] = 32'b00000000011100000100000110000100;
   assign mem[51903:51872] = 32'b11111000000101000010110111101000;
   assign mem[51935:51904] = 32'b00000001011101110010000011010000;
   assign mem[51967:51936] = 32'b00000011001100001011010000001000;
   assign mem[51999:51968] = 32'b11101011111011101001001011000000;
   assign mem[52031:52000] = 32'b00000101100111001010001011001000;
   assign mem[52063:52032] = 32'b11111111011111110001101011001100;
   assign mem[52095:52064] = 32'b00000010011101001001000100001100;
   assign mem[52127:52096] = 32'b00000010110000010001110100110100;
   assign mem[52159:52128] = 32'b00000010101101011100111000001100;
   assign mem[52191:52160] = 32'b00000011111110010010001111110100;
   assign mem[52223:52192] = 32'b00001011111101001000100101110000;
   assign mem[52255:52224] = 32'b11111000100010011100110110100000;
   assign mem[52287:52256] = 32'b11110010110100111001100111100000;
   assign mem[52319:52288] = 32'b00000001100001100100001100100100;
   assign mem[52351:52320] = 32'b11111111111110101011101010010110;
   assign mem[52383:52352] = 32'b00001111010111110111101001110000;
   assign mem[52415:52384] = 32'b11110000111110011011100100010000;
   assign mem[52447:52416] = 32'b11111011111001001001000000101000;
   assign mem[52479:52448] = 32'b11111110101010110000000010011100;
   assign mem[52511:52480] = 32'b00000011000111000011011010000100;
   assign mem[52543:52512] = 32'b11110110011111101110001001000000;
   assign mem[52575:52544] = 32'b00000001101000010110011010001100;
   assign mem[52607:52576] = 32'b00000101101000100000100101011000;
   assign mem[52639:52608] = 32'b11111101111010111001010010110100;
   assign mem[52671:52640] = 32'b11111111100001110011101010001101;
   assign mem[52703:52672] = 32'b11110010110001010010100111100000;
   assign mem[52735:52704] = 32'b00000111011111110011100101101000;
   assign mem[52767:52736] = 32'b00000011001110000000110110001000;
   assign mem[52799:52768] = 32'b00000001011010100011001110011000;
   assign mem[52831:52800] = 32'b00000010001011010100000101010000;
   assign mem[52863:52832] = 32'b11111110110111100111101101000110;
   assign mem[52895:52864] = 32'b11111111011110001010110011100100;
   assign mem[52927:52896] = 32'b00000010001100100100010110000000;
   assign mem[52959:52928] = 32'b00000010100000100111000101011000;
   assign mem[52991:52960] = 32'b11111100000111111101010101101100;
   assign mem[53023:52992] = 32'b11111100010101110010101011000100;
   assign mem[53055:53024] = 32'b11111110100010011111101000101010;
   assign mem[53087:53056] = 32'b11111111101100100111110101011011;
   assign mem[53119:53088] = 32'b11111101001000000001010111111100;
   assign mem[53151:53120] = 32'b11111110011111001111011101100000;
   assign mem[53183:53152] = 32'b00000110000100111111110101110000;
   assign mem[53215:53184] = 32'b00000000101010011000001010001100;
   assign mem[53247:53216] = 32'b00000011110000111011100100010100;
   assign mem[53279:53248] = 32'b11111001001011011000110101111000;
   assign mem[53311:53280] = 32'b00001000010100011010111111000000;
   assign mem[53343:53312] = 32'b11111100001101011001001000110000;
   assign mem[53375:53344] = 32'b00000100110001100000110100110000;
   assign mem[53407:53376] = 32'b11111111011110110100100110111100;
   assign mem[53439:53408] = 32'b11110111100100001101110011010000;
   assign mem[53471:53440] = 32'b11111111110010100010101001110000;
   assign mem[53503:53472] = 32'b11111111001000100111101010011111;
   assign mem[53535:53504] = 32'b11111110000110111101101001011000;
   assign mem[53567:53536] = 32'b00000010001111010001110100001100;
   assign mem[53599:53568] = 32'b11111110111000000100100100101010;
   assign mem[53631:53600] = 32'b11111110100111001101010110100100;
   assign mem[53663:53632] = 32'b11111100010100010010100010111000;
   assign mem[53695:53664] = 32'b11111111000100000000101101111111;
   assign mem[53727:53696] = 32'b00000000101101101011111111000011;
   assign mem[53759:53728] = 32'b00000001100111010111010110011110;
   assign mem[53791:53760] = 32'b11111010100101110111011110111000;
   assign mem[53823:53792] = 32'b11110111010110001001011101110000;
   assign mem[53855:53824] = 32'b00001100011100011100001011000000;
   assign mem[53887:53856] = 32'b00000000000110110001001000010001;
   assign mem[53919:53888] = 32'b11110110110111010110110000100000;
   assign mem[53951:53920] = 32'b00000001111101010111100101100110;
   assign mem[53983:53952] = 32'b11111011011100011011010111101000;
   assign mem[54015:53984] = 32'b11111001011101000000100000111000;
   assign mem[54047:54016] = 32'b11111100000010100011111101011100;
   assign mem[54079:54048] = 32'b11111111011111001100111001101101;
   assign mem[54111:54080] = 32'b11111110101011100011011011011000;
   assign mem[54143:54112] = 32'b00000001001101111110000111111100;
   assign mem[54175:54144] = 32'b11111101011011111101110001110000;
   assign mem[54207:54176] = 32'b00000001110000110100001100010110;
   assign mem[54239:54208] = 32'b11111101000101000111110010101100;
   assign mem[54271:54240] = 32'b00000111001010000010110001110000;
   assign mem[54303:54272] = 32'b00000010011000100111000100110000;
   assign mem[54335:54304] = 32'b11110111111110011001000001000000;
   assign mem[54367:54336] = 32'b00000000011101111010010000100001;
   assign mem[54399:54368] = 32'b11111100000110111011110101110000;
   assign mem[54431:54400] = 32'b11111110011111000010011100001000;
   assign mem[54463:54432] = 32'b11111000111110101011101110100000;
   assign mem[54495:54464] = 32'b00000101100100001001111110111000;
   assign mem[54527:54496] = 32'b00001010010101110000010100000000;
   assign mem[54559:54528] = 32'b11111000000110001100001110110000;
   assign mem[54591:54560] = 32'b11110110011001000101110101110000;
   assign mem[54623:54592] = 32'b11101110011010110010001100000000;
   assign mem[54655:54624] = 32'b00010000101011011101001110100000;
   assign mem[54687:54656] = 32'b00000110100001011110101000010000;
   assign mem[54719:54688] = 32'b11101100000011110110010011000000;
   assign mem[54751:54720] = 32'b11111111001011010001011000001001;
   assign mem[54783:54752] = 32'b00001011000100001010110000100000;
   assign mem[54815:54784] = 32'b11111111001011100101010000011010;
   assign mem[54847:54816] = 32'b00000000000110111001101010001001;
   assign mem[54879:54848] = 32'b00001100000100000001011100100000;
   assign mem[54911:54880] = 32'b11111010011110001010110100111000;
   assign mem[54943:54912] = 32'b00000011111010111110001100110100;
   assign mem[54975:54944] = 32'b00000000011011111111010001111001;
   assign mem[55007:54976] = 32'b11111100001000110000001001011100;
   assign mem[55039:55008] = 32'b11101010100001100001111001100000;
   assign mem[55071:55040] = 32'b11111110111000111001011110100010;
   assign mem[55103:55072] = 32'b00000011010110100110111010110000;
   assign mem[55135:55104] = 32'b11110101010101000101001000110000;
   assign mem[55167:55136] = 32'b00000000101001001111001110001010;
   assign mem[55199:55168] = 32'b11111100101111100011000100010100;
   assign mem[55231:55200] = 32'b00001010101001111000001000110000;
   assign mem[55263:55232] = 32'b11111010111000111000110100111000;
   assign mem[55295:55264] = 32'b11111111110100111010001100110000;
   assign mem[55327:55296] = 32'b00000111000100011000100110001000;
   assign mem[55359:55328] = 32'b11111010111000001100111000101000;
   assign mem[55391:55360] = 32'b11111101110110100101101100001000;
   assign mem[55423:55392] = 32'b00000000001111000110011100101101;
   assign mem[55455:55424] = 32'b00000101001110010110110000111000;
   assign mem[55487:55456] = 32'b00000100000111100101001011110000;
   assign mem[55519:55488] = 32'b00000100011100111001111110111000;
   assign mem[55551:55520] = 32'b11110000110010111000110101000000;
   assign mem[55583:55552] = 32'b11111111000001100100100111111000;
   assign mem[55615:55584] = 32'b11111001111110110101000010110000;
   assign mem[55647:55616] = 32'b00000000000101011010101111111110;
   assign mem[55679:55648] = 32'b00000100101110111110111000100000;
   assign mem[55711:55680] = 32'b11110010111011100110111010100000;
   assign mem[55743:55712] = 32'b00000011000110010001110001001100;
   assign mem[55775:55744] = 32'b00001010010100101000000111110000;
   assign mem[55807:55776] = 32'b00000001011110011000010001101110;
   assign mem[55839:55808] = 32'b00000111001110000100000111101000;
   assign mem[55871:55840] = 32'b11111011111010100111011001111000;
   assign mem[55903:55872] = 32'b11111110101110011001110010100100;
   assign mem[55935:55904] = 32'b11100000101001011001010001000000;
   assign mem[55967:55936] = 32'b00000001100111010011100111100110;
   assign mem[55999:55968] = 32'b11100110000001101010000001100000;
   assign mem[56031:56000] = 32'b11111100011111110111001010101000;
   assign mem[56063:56032] = 32'b11111100011110010010010110010000;
   assign mem[56095:56064] = 32'b00000001111110010011100111111010;
   assign mem[56127:56096] = 32'b11111101100000001101101101110100;
   assign mem[56159:56128] = 32'b11111111110001100001101001111000;
   assign mem[56191:56160] = 32'b11111101001101010001110110000100;
   assign mem[56223:56192] = 32'b11111110110101100100111001111010;
   assign mem[56255:56224] = 32'b00000010110001010000111000000100;
   assign mem[56287:56256] = 32'b00000000010101110111011010110101;
   assign mem[56319:56288] = 32'b11111101010010010000100110010000;
   assign mem[56351:56320] = 32'b00000110110010000101111110110000;
   assign mem[56383:56352] = 32'b11111001001000111011001010100000;
   assign mem[56415:56384] = 32'b00000111100111110000100110110000;
   assign mem[56447:56416] = 32'b11111011011100001111011100110000;
   assign mem[56479:56448] = 32'b11110010101001010110000100010000;
   assign mem[56511:56480] = 32'b00000111001010001100110010011000;
   assign mem[56543:56512] = 32'b11111000011010001011010000001000;
   assign mem[56575:56544] = 32'b00000000100000010110000111001100;
   assign mem[56607:56576] = 32'b00000000001010100000011001000110;
   assign mem[56639:56608] = 32'b00000010001010001100011001010100;
   assign mem[56671:56640] = 32'b11111111100110011001111001011110;
   assign mem[56703:56672] = 32'b11111110110110111101010101011110;
   assign mem[56735:56704] = 32'b11111111110101011001101110001111;
   assign mem[56767:56736] = 32'b11111001110011010000000110110000;
   assign mem[56799:56768] = 32'b11111110111100101000010001100110;
   assign mem[56831:56800] = 32'b11111110001010100111000010100100;
   assign mem[56863:56832] = 32'b11111101111111000000111001010100;
   assign mem[56895:56864] = 32'b11111100000110011111101000011000;
   assign mem[56927:56896] = 32'b00000000001011000001000100000100;
   assign mem[56959:56928] = 32'b00000000111011011101010101111011;
   assign mem[56991:56960] = 32'b00000000011100110001010000100111;
   assign mem[57023:56992] = 32'b00000101001001101000010011000000;
   assign mem[57055:57024] = 32'b00000110101000011010100011111000;
   assign mem[57087:57056] = 32'b11111111010111101011010101001001;
   assign mem[57119:57088] = 32'b11111110001100010011111111010110;
   assign mem[57151:57120] = 32'b11111101110101110110011011000100;
   assign mem[57183:57152] = 32'b11111111101110110100001010010011;
   assign mem[57215:57184] = 32'b11110110101000000110001001100000;
   assign mem[57247:57216] = 32'b00000000111010101101011101111010;
   assign mem[57279:57248] = 32'b00000001010010111100010101101100;
   assign mem[57311:57280] = 32'b00000010111100001001010101100100;
   assign mem[57343:57312] = 32'b00000110001010010001100100011000;
   assign mem[57375:57344] = 32'b11111100100110001011000111001000;
   assign mem[57407:57376] = 32'b00000101010001000001011001111000;
   assign mem[57439:57408] = 32'b00000001111111011100001000001100;
   assign mem[57471:57440] = 32'b11111101011101110000101001111000;
   assign mem[57503:57472] = 32'b00000010011010110101000011111000;
   assign mem[57535:57504] = 32'b11110010101001011101111001000000;
   assign mem[57567:57536] = 32'b11111110000010000100101110000100;
   assign mem[57599:57568] = 32'b11111001000111001101011111101000;
   assign mem[57631:57600] = 32'b11111110001100000100101101010010;
   assign mem[57663:57632] = 32'b11111010011001000000010101101000;
   assign mem[57695:57664] = 32'b11111110100010001100101010100100;
   assign mem[57727:57696] = 32'b00000111101010110001011101110000;
   assign mem[57759:57728] = 32'b11101110011110111110010011100000;
   assign mem[57791:57760] = 32'b00000100111111110000001011101000;
   assign mem[57823:57792] = 32'b00000000001100101100101100001111;
   assign mem[57855:57824] = 32'b00000100110000011111011101000000;
   assign mem[57887:57856] = 32'b00000000101000011000111000000010;
   assign mem[57919:57888] = 32'b00000001000001110000110001111000;
   assign mem[57951:57920] = 32'b11111101000000100101010111001100;
   assign mem[57983:57952] = 32'b11110111100001011001110111010000;
   assign mem[58015:57984] = 32'b00000000010001001111100100000110;
   assign mem[58047:58016] = 32'b00000100110010000001101101010000;
   assign mem[58079:58048] = 32'b11110111101101111001101000000000;
   assign mem[58111:58080] = 32'b00000100000101110100111110101000;
   assign mem[58143:58112] = 32'b11110110111000011010110110100000;
   assign mem[58175:58144] = 32'b00000100001111011011111110010000;
   assign mem[58207:58176] = 32'b00000001001110011100111010011110;
   assign mem[58239:58208] = 32'b00000100011010011000001101010000;
   assign mem[58271:58240] = 32'b00000100000010001100001101110000;
   assign mem[58303:58272] = 32'b11111110000110000011000010101110;
   assign mem[58335:58304] = 32'b00000101000001011111000110100000;
   assign mem[58367:58336] = 32'b11111111011111111011011111101101;
   assign mem[58399:58368] = 32'b11100110100010011010001010000000;
   assign mem[58431:58400] = 32'b00000101101111111010001100000000;
   assign mem[58463:58432] = 32'b00000000100101101111111110101001;
   assign mem[58495:58464] = 32'b00000000111101110011010101011010;
   assign mem[58527:58496] = 32'b11111100100110110010100011010100;
   assign mem[58559:58528] = 32'b00000100100101000100110111111000;
   assign mem[58591:58560] = 32'b11111100101111011100111001001000;
   assign mem[58623:58592] = 32'b00001001010100011000010000010000;
   assign mem[58655:58624] = 32'b11110011111101001110000000110000;
   assign mem[58687:58656] = 32'b11110000011100001111010000000000;
   assign mem[58719:58688] = 32'b00010011100001011011011101100000;
   assign mem[58751:58720] = 32'b11111100100111011001001101110000;
   assign mem[58783:58752] = 32'b00001101110011000001100011000000;
   assign mem[58815:58784] = 32'b11100100011011110011001111000000;
   assign mem[58847:58816] = 32'b11111111000101110100000001111001;
   assign mem[58879:58848] = 32'b11101101101010101111001011100000;
   assign mem[58911:58880] = 32'b11111010101101101011100111000000;
   assign mem[58943:58912] = 32'b00000101100001000010111111110000;
   assign mem[58975:58944] = 32'b11111111001100000101010100010000;
   assign mem[59007:58976] = 32'b00001011000011010110100001100000;
   assign mem[59039:59008] = 32'b11111101110111011000011011101000;
   assign mem[59071:59040] = 32'b11111000111000000011011110011000;
   assign mem[59103:59072] = 32'b00001000100011010111010010110000;
   assign mem[59135:59104] = 32'b11110001101101010011100100100000;
   assign mem[59167:59136] = 32'b00000100101000101011001110010000;
   assign mem[59199:59168] = 32'b11110000101101000000010110110000;
   assign mem[59231:59200] = 32'b11111000010011011100101001001000;
   assign mem[59263:59232] = 32'b00000001010001001110001111011010;
   assign mem[59295:59264] = 32'b00000011100100111110111101110100;
   assign mem[59327:59296] = 32'b00001010100010001100101010000000;
   assign mem[59359:59328] = 32'b00000000111110100110000001001100;
   assign mem[59391:59360] = 32'b11110101111100100001001011000000;
   assign mem[59423:59392] = 32'b11111100001101001110110111001100;
   assign mem[59455:59424] = 32'b11111111010011100100100101101010;
   assign mem[59487:59456] = 32'b00000011111100001110010010000000;
   assign mem[59519:59488] = 32'b11101000011011010100110111000000;
   assign mem[59551:59520] = 32'b00000011110000101001100010011100;
   assign mem[59583:59552] = 32'b00000100000011100000111110100000;
   assign mem[59615:59584] = 32'b11111111011000101010000010101110;
   assign mem[59647:59616] = 32'b00000000110000011011010010101111;
   assign mem[59679:59648] = 32'b00000010011111100111111100111000;
   assign mem[59711:59680] = 32'b11111111011011000111001101110110;
   assign mem[59743:59712] = 32'b11111110010001111101001110101000;
   assign mem[59775:59744] = 32'b00000000101101001000100010001000;
   assign mem[59807:59776] = 32'b11111100101010001110110100000000;
   assign mem[59839:59808] = 32'b00000000001010110011001001110010;
   assign mem[59871:59840] = 32'b00000010000011110101000001011000;
   assign mem[59903:59872] = 32'b00000100011100000111010101110000;
   assign mem[59935:59904] = 32'b00000101000100111011101011000000;
   assign mem[59967:59936] = 32'b00000011000001111101111011100000;
   assign mem[59999:59968] = 32'b00000000000110100101011100111000;
   assign mem[60031:60000] = 32'b11111101010010101010010101110100;
   assign mem[60063:60032] = 32'b11111100000010111011011011100000;
   assign mem[60095:60064] = 32'b00000000100100001000100010100110;
   assign mem[60127:60096] = 32'b00000000101111100111001101011000;
   assign mem[60159:60128] = 32'b00000011110100110110111000010000;
   assign mem[60191:60160] = 32'b11111111110111001011111011010000;
   assign mem[60223:60192] = 32'b00000001111001101001001100011110;
   assign mem[60255:60224] = 32'b00000000111101000011001100001001;
   assign mem[60287:60256] = 32'b11111110000010110001100101111000;
   assign mem[60319:60288] = 32'b00000000101010011101001101100101;
   assign mem[60351:60320] = 32'b11111110111011111001110000001000;
   assign mem[60383:60352] = 32'b11111010101000011101111000001000;
   assign mem[60415:60384] = 32'b00000010010110011101100111000000;
   assign mem[60447:60416] = 32'b00000010000010010010111110100100;
   assign mem[60479:60448] = 32'b00000010111000001001100010110000;
   assign mem[60511:60480] = 32'b11111101100000000000100100110000;
   assign mem[60543:60512] = 32'b00000000011111100110001010110111;
   assign mem[60575:60544] = 32'b00000001100111001110101011000100;
   assign mem[60607:60576] = 32'b11111000110011111101100001110000;
   assign mem[60639:60608] = 32'b00000000011001000010011111001111;
   assign mem[60671:60640] = 32'b11111110011101100000001000010110;
   assign mem[60703:60672] = 32'b00000100100100011011110100000000;
   assign mem[60735:60704] = 32'b11111001001111101101111010110000;
   assign mem[60767:60736] = 32'b00000000000101000100010010110111;
   assign mem[60799:60768] = 32'b00000011100111100101001110011000;
   assign mem[60831:60800] = 32'b00000000010100111000010101011100;
   assign mem[60863:60832] = 32'b00000110010011000010011001110000;
   assign mem[60895:60864] = 32'b11111100101001010011010001010000;
   assign mem[60927:60896] = 32'b11111010111001110011100011000000;
   assign mem[60959:60928] = 32'b00000100100001001101000001100000;
   assign mem[60991:60960] = 32'b00000011100001100000000001100100;
   assign mem[61023:60992] = 32'b00000110100101101001101110110000;
   assign mem[61055:61024] = 32'b11110011011100011111111010000000;
   assign mem[61087:61056] = 32'b11111001101100110101100000000000;
   assign mem[61119:61088] = 32'b11111111000011000110111111011010;
   assign mem[61151:61120] = 32'b00000000100101100111011110011100;
   assign mem[61183:61152] = 32'b00000111011010100010110101111000;
   assign mem[61215:61184] = 32'b11111001100110100101000110001000;
   assign mem[61247:61216] = 32'b11111010101011110111100101001000;
   assign mem[61279:61248] = 32'b00001000001000111011001100000000;
   assign mem[61311:61280] = 32'b00000110001000100011011000101000;
   assign mem[61343:61312] = 32'b00000010111101101011000010100100;
   assign mem[61375:61344] = 32'b00000000101101000000111101011111;
   assign mem[61407:61376] = 32'b11111010111111101001100010110000;
   assign mem[61439:61408] = 32'b11110111001110101101100000110000;
   assign mem[61471:61440] = 32'b11111111100100101001100100000000;
   assign mem[61503:61472] = 32'b11111010101011101000111001001000;
   assign mem[61535:61504] = 32'b11111110011011010111111101101010;
   assign mem[61567:61536] = 32'b00000110011111111100001011011000;
   assign mem[61599:61568] = 32'b11111110000100000001101100100010;
   assign mem[61631:61600] = 32'b11111111100110011001110110000010;
   assign mem[61663:61632] = 32'b11111010010101101101110011001000;
   assign mem[61695:61664] = 32'b00000011011101001010010010101000;
   assign mem[61727:61696] = 32'b00000001001100010111001000101100;
   assign mem[61759:61728] = 32'b00000001110010100110110000101100;
   assign mem[61791:61760] = 32'b00000001011011000101010001010110;
   assign mem[61823:61792] = 32'b00000000101100001110110100111010;
   assign mem[61855:61824] = 32'b00000001001110111000001001011010;
   assign mem[61887:61856] = 32'b00000001101110100111001010111100;
   assign mem[61919:61888] = 32'b00000100011101111001111111101000;
   assign mem[61951:61920] = 32'b11111010010010110100111101100000;
   assign mem[61983:61952] = 32'b11111010011011011101101100000000;
   assign mem[62015:61984] = 32'b11111101110100000111011000000100;
   assign mem[62047:62016] = 32'b00000001010101000011110011000000;
   assign mem[62079:62048] = 32'b00000000010010100110110000010111;
   assign mem[62111:62080] = 32'b00000101111100001101000011010000;
   assign mem[62143:62112] = 32'b11110100011100000110000110010000;
   assign mem[62175:62144] = 32'b00000100101110010111111100100000;
   assign mem[62207:62176] = 32'b00000101100010011100010101000000;
   assign mem[62239:62208] = 32'b11110010011011011000101110100000;
   assign mem[62271:62240] = 32'b11111110110100010110001100101010;
   assign mem[62303:62272] = 32'b11111110101011011000010110101110;
   assign mem[62335:62304] = 32'b00000001000011111111001011001110;
   assign mem[62367:62336] = 32'b00000010000110110101111000001000;
   assign mem[62399:62368] = 32'b00000001010010111101001110110000;
   assign mem[62431:62400] = 32'b11111110111011000101111000110010;
   assign mem[62463:62432] = 32'b00000010011110101011010110010000;
   assign mem[62495:62464] = 32'b11111011110011001101101100101000;
   assign mem[62527:62496] = 32'b00000110000101110101001010101000;
   assign mem[62559:62528] = 32'b11111000111011000110010111100000;
   assign mem[62591:62560] = 32'b00000001101011001110101011000000;
   assign mem[62623:62592] = 32'b11111011100110111101101011110000;
   assign mem[62655:62624] = 32'b11111011000010100101010001000000;
   assign mem[62687:62656] = 32'b11111010110001011110001011011000;
   assign mem[62719:62688] = 32'b11111110111010100011000110100000;
   assign mem[62751:62720] = 32'b11111101110001000000000000000100;
   assign mem[62783:62752] = 32'b00001001111001111101100100100000;
   assign mem[62815:62784] = 32'b11111001110001111010111111000000;
   assign mem[62847:62816] = 32'b11110011110011010010101111000000;
   assign mem[62879:62848] = 32'b11111010111100011011111111000000;
   assign mem[62911:62880] = 32'b00001110000111111110011011100000;
   assign mem[62943:62912] = 32'b00000110010110111011110001011000;
   assign mem[62975:62944] = 32'b11111110001101101111001100110110;
   assign mem[63007:62976] = 32'b11111010101010000100011001101000;
   assign mem[63039:63008] = 32'b11100110111100000001011111000000;
   assign mem[63071:63040] = 32'b00000000000010010010101001100111;
   assign mem[63103:63072] = 32'b00000011000010111011101101101100;
   assign mem[63135:63104] = 32'b00000001010001100100001000101110;
   assign mem[63167:63136] = 32'b11110111111010011111011000010000;
   assign mem[63199:63168] = 32'b11111000111001101100011000010000;
   assign mem[63231:63200] = 32'b11111101010101110010101011110100;
   assign mem[63263:63232] = 32'b00000100010101111101001001101000;
   assign mem[63295:63264] = 32'b11111001011110100101010100001000;
   assign mem[63327:63296] = 32'b00000010100000000101011100010000;
   assign mem[63359:63328] = 32'b11111001111000111001100110101000;
   assign mem[63391:63360] = 32'b11110111001000100010010001110000;
   assign mem[63423:63392] = 32'b00001010110110011101000011000000;
   assign mem[63455:63424] = 32'b11110100100000101011110000100000;
   assign mem[63487:63456] = 32'b00000100111111010011100011000000;
   assign mem[63519:63488] = 32'b00000101000100100101101000110000;
   assign mem[63551:63520] = 32'b11111001100111101010111100010000;
   assign mem[63583:63552] = 32'b00000110011010010111111101011000;
   assign mem[63615:63584] = 32'b11111011101111110010110001110000;
   assign mem[63647:63616] = 32'b11111001001010100101111001001000;
   assign mem[63679:63648] = 32'b11110001011000100101100001110000;
   assign mem[63711:63680] = 32'b11110110110001001010111011110000;
   assign mem[63743:63712] = 32'b00001000000111101011110000010000;
   assign mem[63775:63744] = 32'b11110001100010101011101100100000;
   assign mem[63807:63776] = 32'b11110010111010111101110000100000;
   assign mem[63839:63808] = 32'b00000111110100111010001101111000;
   assign mem[63871:63840] = 32'b11111111111111000101101101000100;
   assign mem[63903:63872] = 32'b00000101101001100101110001001000;
   assign mem[63935:63904] = 32'b00000000001101011010000100110000;
   assign mem[63967:63936] = 32'b11111111110000010101111111111100;
   assign mem[63999:63968] = 32'b11110110101001000111111010010000;
   assign mem[64031:64000] = 32'b00000001100001110111010100000010;
   assign mem[64063:64032] = 32'b00000010000000000011000101010000;
   assign mem[64095:64064] = 32'b11111111010111000100101110111101;
   assign mem[64127:64096] = 32'b00000001010011101111011101000000;
   assign mem[64159:64128] = 32'b00000001001010100111100010000010;
   assign mem[64191:64160] = 32'b11111110011010100100000011010000;
   assign mem[64223:64192] = 32'b11111011010001100000001010011000;
   assign mem[64255:64224] = 32'b00000001010100111010001110111100;
   assign mem[64287:64256] = 32'b00000001101010000111100000101010;
   assign mem[64319:64288] = 32'b00000001111110011101100001010100;
   assign mem[64351:64320] = 32'b11111011101111011011001001110000;
   assign mem[64383:64352] = 32'b00010001111111001010011111100000;
   assign mem[64415:64384] = 32'b11110010001111010011111111110000;
   assign mem[64447:64416] = 32'b11111011010001101011000110011000;
   assign mem[64479:64448] = 32'b00001010110110100010101011110000;
   assign mem[64511:64480] = 32'b00000000101010010011000010000111;
   assign mem[64543:64512] = 32'b00000010100100110000011111000100;
   assign mem[64575:64544] = 32'b11101101001100110010000100000000;
   assign mem[64607:64576] = 32'b11111111110111100110111011001101;
   assign mem[64639:64608] = 32'b11110011000001101001011101100000;
   assign mem[64671:64640] = 32'b11111010101001101011010010011000;
   assign mem[64703:64672] = 32'b11111100001101011111110111110000;
   assign mem[64735:64704] = 32'b00000010111000000001101111011100;
   assign mem[64767:64736] = 32'b11111110111101001100111010011100;
   assign mem[64799:64768] = 32'b11110111001010110100101110100000;
   assign mem[64831:64800] = 32'b00000010110010111111110111110100;
   assign mem[64863:64832] = 32'b11111101101110111111100101100000;
   assign mem[64895:64864] = 32'b11111111110010000111101111101000;
   assign mem[64927:64896] = 32'b00000001001100110001100001000000;
   assign mem[64959:64928] = 32'b00000010111001011010101111101100;
   assign mem[64991:64960] = 32'b11111101000100000100100101010000;
   assign mem[65023:64992] = 32'b11111001010110100111011001110000;
   assign mem[65055:65024] = 32'b11111111111011001010101101100001;
   assign mem[65087:65056] = 32'b00000001010001111101001011111100;
   assign mem[65119:65088] = 32'b00000001001100110100000111100100;
   assign mem[65151:65120] = 32'b11111011100101101000100010101000;
   assign mem[65183:65152] = 32'b11111110100100110011011011111100;
   assign mem[65215:65184] = 32'b11111111011101011000000100011010;
   assign mem[65247:65216] = 32'b11111111000010011110011000010101;
   assign mem[65279:65248] = 32'b00000010001111111001011011110000;
   assign mem[65311:65280] = 32'b11111011110101010101110001011000;
   assign mem[65343:65312] = 32'b11111011100011000011010101001000;
   assign mem[65375:65344] = 32'b00000000001001110111001100000110;
   assign mem[65407:65376] = 32'b00000110000000010000010111000000;
   assign mem[65439:65408] = 32'b11111000101111110010001010010000;
   assign mem[65471:65440] = 32'b00000011100011110001110101101100;
   assign mem[65503:65472] = 32'b11111001010101000110011101010000;
   assign mem[65535:65504] = 32'b00000010110001000110111101001000;
   assign mem[65567:65536] = 32'b00000000011110111100100110101111;
   assign mem[65599:65568] = 32'b00000011100100011100000111100000;
   assign mem[65631:65600] = 32'b11111101100000011101100010100100;
   assign mem[65663:65632] = 32'b11111110001000011001000001010110;
   assign mem[65695:65664] = 32'b11111110101101100100000101000110;
   assign mem[65727:65696] = 32'b00000001100001001100000000011000;
   assign mem[65759:65728] = 32'b11111101001010111001110100001000;
   assign mem[65791:65760] = 32'b00000010011011110000110000000100;
   assign mem[65823:65792] = 32'b11111101011111110110100001010000;
   assign mem[65855:65824] = 32'b00000000111000010001010110101111;
   assign mem[65887:65856] = 32'b00000000001011000001000111011111;
   assign mem[65919:65888] = 32'b00000100010100001101101100010000;
   assign mem[65951:65920] = 32'b00000011010000001111101010010100;
   assign mem[65983:65952] = 32'b11111101110100100100100100011100;
   assign mem[66015:65984] = 32'b11111101110010000011010000101000;
   assign mem[66047:66016] = 32'b00000011011000100000000111010100;
   assign mem[66079:66048] = 32'b11101110100101011111000101100000;
   assign mem[66111:66080] = 32'b00000000100011110011111110011000;
   assign mem[66143:66112] = 32'b11111101011000010010011000011000;
   assign mem[66175:66144] = 32'b00000111000110001100110110000000;
   assign mem[66207:66176] = 32'b11111100101100101110000111000100;
   assign mem[66239:66208] = 32'b00000010100000110011011111011000;
   assign mem[66271:66240] = 32'b11111101000111100001101111001100;
   assign mem[66303:66272] = 32'b00000101000010001110101110100000;
   assign mem[66335:66304] = 32'b11111010111100010010110001110000;
   assign mem[66367:66336] = 32'b11101101011101100011100010000000;
   assign mem[66399:66368] = 32'b00001001101000000110101100010000;
   assign mem[66431:66400] = 32'b11111111111011110010111100000110;
   assign mem[66463:66432] = 32'b00000101111010101101101011101000;
   assign mem[66495:66464] = 32'b11110111101001110010111001000000;
   assign mem[66527:66496] = 32'b00000010010000111001010011010000;
   assign mem[66559:66528] = 32'b11111000110101100000010100111000;
   assign mem[66591:66560] = 32'b11111101111110011100000010000100;
   assign mem[66623:66592] = 32'b00000000110010111110100000000001;
   assign mem[66655:66624] = 32'b11111100110011111000001101100100;
   assign mem[66687:66656] = 32'b11111101111011110111011001101000;
   assign mem[66719:66688] = 32'b11111010101010100001000111010000;
   assign mem[66751:66720] = 32'b00001011001010110001011100010000;
   assign mem[66783:66752] = 32'b11111100011111010100011100000000;
   assign mem[66815:66784] = 32'b11111101000100010111010100111100;
   assign mem[66847:66816] = 32'b11111100100101100111111110101000;
   assign mem[66879:66848] = 32'b11111101101000010110111101010100;
   assign mem[66911:66880] = 32'b00000000101110101111011011000010;
   assign mem[66943:66912] = 32'b11111011110010100110110011011000;
   assign mem[66975:66944] = 32'b00000011011111101001110011011100;
   assign mem[67007:66976] = 32'b00000110110011011000001001010000;
   assign mem[67039:67008] = 32'b11101001111100100001110010000000;
   assign mem[67071:67040] = 32'b11111111011011110110000111110101;
   assign mem[67103:67072] = 32'b11111101111011001010000110110100;
   assign mem[67135:67104] = 32'b11111110111100100111011010100100;
   assign mem[67167:67136] = 32'b00000010101000110001011100011000;
   assign mem[67199:67168] = 32'b00000000111011010110000010110000;
   assign mem[67231:67200] = 32'b00000000111001110111001001001101;
   assign mem[67263:67232] = 32'b00000001100101101110111100101010;
   assign mem[67295:67264] = 32'b00000011101010111011000111110000;
   assign mem[67327:67296] = 32'b11111111010011000001000100011111;
   assign mem[67359:67328] = 32'b00000000010100011000100101101100;
   assign mem[67391:67360] = 32'b11110110101011001101111000000000;
   assign mem[67423:67392] = 32'b11111011001100101000011001000000;
   assign mem[67455:67424] = 32'b11111111101010001110101101010000;
   assign mem[67487:67456] = 32'b11111010011000101111110001110000;
   assign mem[67519:67488] = 32'b00000010101100011100100011110000;
   assign mem[67551:67520] = 32'b11111111100101001001010110101001;
   assign mem[67583:67552] = 32'b11111101111100001101110111111100;
   assign mem[67615:67584] = 32'b00000011100000110101100111100100;
   assign mem[67647:67616] = 32'b11111111011110010111001111001001;
   assign mem[67679:67648] = 32'b11111100000010111000111101111100;
   assign mem[67711:67680] = 32'b00000010011000101000101011010000;
   assign mem[67743:67712] = 32'b11111011010011111100110101010000;
   assign mem[67775:67744] = 32'b00000000111100110100010010111001;
   assign mem[67807:67776] = 32'b11111110111011111110000100011110;
   assign mem[67839:67808] = 32'b00000100110011001110011001011000;
   assign mem[67871:67840] = 32'b11111101010000101011111011001000;
   assign mem[67903:67872] = 32'b00000001010011101011101001011100;
   assign mem[67935:67904] = 32'b00000010110001110110011000001000;
   assign mem[67967:67936] = 32'b11111011011010001001000010110000;
   assign mem[67999:67968] = 32'b00000111010100110111101110101000;
   assign mem[68031:68000] = 32'b00000000101101111101101110101000;
   assign mem[68063:68032] = 32'b00000001111011001111001010001000;
   assign mem[68095:68064] = 32'b11110100001111010000001111000000;
   assign mem[68127:68096] = 32'b00000010011100100101100100011100;
   assign mem[68159:68128] = 32'b11110001110100100001100111000000;
   assign mem[68191:68160] = 32'b00000000001100111010110101011111;
   assign mem[68223:68192] = 32'b11111111101101011111001101000111;
   assign mem[68255:68224] = 32'b00000000010001001011001010100010;
   assign mem[68287:68256] = 32'b11111100011111011010010110101100;
   assign mem[68319:68288] = 32'b11111010110000000001011010101000;
   assign mem[68351:68320] = 32'b00000100000010001010100100101000;
   assign mem[68383:68352] = 32'b00000000100001100101011100010011;
   assign mem[68415:68384] = 32'b00000011001010011010010000110100;
   assign mem[68447:68416] = 32'b11111111010011110100110111111011;
   assign mem[68479:68448] = 32'b00000011000101100010101000011100;
   assign mem[68511:68480] = 32'b11111101000100101110000110010100;
   assign mem[68543:68512] = 32'b00000011000100010001000101011100;
   assign mem[68575:68544] = 32'b11110110000001111010100010000000;
   assign mem[68607:68576] = 32'b11111001100111100100000011100000;
   assign mem[68639:68608] = 32'b00001000101111101011010111010000;
   assign mem[68671:68640] = 32'b11111011110000111100110100111000;
   assign mem[68703:68672] = 32'b00000111011010000110001111000000;
   assign mem[68735:68704] = 32'b00000110000000001000111111101000;
   assign mem[68767:68736] = 32'b11111101111111101000011110100000;
   assign mem[68799:68768] = 32'b11111001000001001011110010001000;
   assign mem[68831:68800] = 32'b00000111100110010110111000001000;
   assign mem[68863:68832] = 32'b11111101000111000011001100010000;
   assign mem[68895:68864] = 32'b00000111111101010011011100010000;
   assign mem[68927:68896] = 32'b00000010000000101101010010110000;
   assign mem[68959:68928] = 32'b00000110111100101111010110101000;
   assign mem[68991:68960] = 32'b11110111100000001101100010100000;
   assign mem[69023:68992] = 32'b11111010000001001010111011011000;
   assign mem[69055:69024] = 32'b11111111001101000011011000010011;
   assign mem[69087:69056] = 32'b11111100010001011111001100100100;
   assign mem[69119:69088] = 32'b11111100001110001111100100110100;
   assign mem[69151:69120] = 32'b00000100011111100111101000110000;
   assign mem[69183:69152] = 32'b00000001100101111100001001111000;
   assign mem[69215:69184] = 32'b00000100011111101100111011010000;
   assign mem[69247:69216] = 32'b00000010111010000100010001001000;
   assign mem[69279:69248] = 32'b00001100110000100101100011100000;
   assign mem[69311:69280] = 32'b11110111110101111100101111010000;
   assign mem[69343:69312] = 32'b11111110000001110101011111111010;
   assign mem[69375:69344] = 32'b11111000011111110110100101000000;
   assign mem[69407:69376] = 32'b00000010101011010011100010011100;
   assign mem[69439:69408] = 32'b11110000011010100000010010000000;
   assign mem[69471:69440] = 32'b11111101110111010010110001001000;
   assign mem[69503:69472] = 32'b00000111100001001011100000000000;
   assign mem[69535:69504] = 32'b00000110100111100001001110110000;
   assign mem[69567:69536] = 32'b00000110001000100111001010011000;
   assign mem[69599:69568] = 32'b11111101001101110111100101101000;
   assign mem[69631:69600] = 32'b11110001101100101001000111010000;
   assign mem[69663:69632] = 32'b00000100000011010001100111101000;
   assign mem[69695:69664] = 32'b11111101001100100111100110101000;
   assign mem[69727:69696] = 32'b11111010001011110010001011100000;
   assign mem[69759:69728] = 32'b11110111001110011001001010010000;
   assign mem[69791:69760] = 32'b11111001010111011010000011000000;
   assign mem[69823:69792] = 32'b00001000011001101110111010010000;
   assign mem[69855:69824] = 32'b00000010110101000101010010111000;
   assign mem[69887:69856] = 32'b11111000011110100100001001110000;
   assign mem[69919:69888] = 32'b00000101101111000110000101111000;
   assign mem[69951:69920] = 32'b11111000010101111010100000111000;
   assign mem[69983:69952] = 32'b11111110101101010101000000100000;
   assign mem[70015:69984] = 32'b11111100000000101011010011001000;
   assign mem[70047:70016] = 32'b11111110110010110000110010110110;
   assign mem[70079:70048] = 32'b11110101111001100110010111100000;
   assign mem[70111:70080] = 32'b00000011001101001000101111100000;
   assign mem[70143:70112] = 32'b00000100111001000001001110110000;
   assign mem[70175:70144] = 32'b11111011011101111111000100101000;
   assign mem[70207:70176] = 32'b11110111111101100010011100010000;
   assign mem[70239:70208] = 32'b00000101111011111001101000011000;
   assign mem[70271:70240] = 32'b00000100100010101101101110111000;
   assign mem[70303:70272] = 32'b00000000110100110000000010001101;
   assign mem[70335:70304] = 32'b11111100100111101110101010100100;
   assign mem[70367:70336] = 32'b00000001111100100110010100100010;
   assign mem[70399:70368] = 32'b00000000100110010100101010000010;
   assign mem[70431:70400] = 32'b11111101110100011001010010010000;
   assign mem[70463:70432] = 32'b11111110001110100011001111010010;
   assign mem[70495:70464] = 32'b11111101101101000110100000010000;
   assign mem[70527:70496] = 32'b00000000111001100001010111001001;
   assign mem[70559:70528] = 32'b11110101011011001001000100100000;
   assign mem[70591:70560] = 32'b00000001110110010001100001000110;
   assign mem[70623:70592] = 32'b11111010000000010100011110001000;
   assign mem[70655:70624] = 32'b00000101001110101001001010110000;
   assign mem[70687:70656] = 32'b00000000001100110010110011001100;
   assign mem[70719:70688] = 32'b00000001110110010101101000111100;
   assign mem[70751:70720] = 32'b11111110011010010100000111011000;
   assign mem[70783:70752] = 32'b11111011010101010111011001010000;
   assign mem[70815:70784] = 32'b11111101010011101110001110001100;
   assign mem[70847:70816] = 32'b00000000100000101010110110010001;
   assign mem[70879:70848] = 32'b11111001100110000000100000101000;
   assign mem[70911:70880] = 32'b11111110111110001000010111011100;
   assign mem[70943:70912] = 32'b11111011000100000110110111010000;
   assign mem[70975:70944] = 32'b00000011000010110000000001101000;
   assign mem[71007:70976] = 32'b00000000011100000111111110000101;
   assign mem[71039:71008] = 32'b00000001011111111110111111101110;
   assign mem[71071:71040] = 32'b11111101011101110000001010101000;
   assign mem[71103:71072] = 32'b00000101001001011101011010001000;
   assign mem[71135:71104] = 32'b00000110011111010000111000001000;
   assign mem[71167:71136] = 32'b11111111010001110001101100000111;
   assign mem[71199:71168] = 32'b00001010001000110100111110110000;
   assign mem[71231:71200] = 32'b11111101001011100111000001011100;
   assign mem[71263:71232] = 32'b00000010101111100110011101101000;
   assign mem[71295:71264] = 32'b00000000000110111011001110010011;
   assign mem[71327:71296] = 32'b11111000101010000000111111110000;
   assign mem[71359:71328] = 32'b11110101111101010010111100010000;
   assign mem[71391:71360] = 32'b11111110101111101010101101001110;
   assign mem[71423:71392] = 32'b11111010011001111001110011011000;
   assign mem[71455:71424] = 32'b11111110110110101101101101011010;
   assign mem[71487:71456] = 32'b11111101110100001110010110010100;
   assign mem[71519:71488] = 32'b11110010010011101111011101110000;
   assign mem[71551:71520] = 32'b00000110111111110111101110111000;
   assign mem[71583:71552] = 32'b00000011011011000100100110011100;
   assign mem[71615:71584] = 32'b00000001001000100001110011010110;
   assign mem[71647:71616] = 32'b11111100011101101000010010101000;
   assign mem[71679:71648] = 32'b00000101100010010010111010010000;
   assign mem[71711:71680] = 32'b00000000100001110000101100010001;
   assign mem[71743:71712] = 32'b00001000111110000111001101100000;
   assign mem[71775:71744] = 32'b11111111000111001111110101001010;
   assign mem[71807:71776] = 32'b00000000110001101101001111101010;
   assign mem[71839:71808] = 32'b11111110000010111011111010000110;
   assign mem[71871:71840] = 32'b00000000010000000001110000100101;
   assign mem[71903:71872] = 32'b00000001111010000100100110011010;
   assign mem[71935:71904] = 32'b00000001010101100001100110000100;
   assign mem[71967:71936] = 32'b11111011100000001110010000011000;
   assign mem[71999:71968] = 32'b00000000101111110100110111111010;
   assign mem[72031:72000] = 32'b00001000001100111111001110110000;
   assign mem[72063:72032] = 32'b00000111111101111101010001100000;
   assign mem[72095:72064] = 32'b11110101110101101011000011110000;
   assign mem[72127:72096] = 32'b11110011101011011010101000110000;
   assign mem[72159:72128] = 32'b00000111000100011100101101111000;
   assign mem[72191:72160] = 32'b00000000001000011110010011011111;
   assign mem[72223:72192] = 32'b00000111011100000011110111000000;
   assign mem[72255:72224] = 32'b11111101111110110011010111001100;
   assign mem[72287:72256] = 32'b00000000101001101000100001000001;
   assign mem[72319:72288] = 32'b11111011000000011011111101010000;
   assign mem[72351:72320] = 32'b11111001011101101110110101000000;
   assign mem[72383:72352] = 32'b11110000101111110101110100010000;
   assign mem[72415:72384] = 32'b00000000001010010010101000100001;
   assign mem[72447:72416] = 32'b00000010000011101100110111100100;
   assign mem[72479:72448] = 32'b11101000011111101000000000000000;
   assign mem[72511:72480] = 32'b00000110011001010011111001111000;
   assign mem[72543:72512] = 32'b00000010110101110111001101011000;
   assign mem[72575:72544] = 32'b11111101011111001100000001101100;
   assign mem[72607:72576] = 32'b00000100110111010101100011100000;
   assign mem[72639:72608] = 32'b00000101000001111110010100101000;
   assign mem[72671:72640] = 32'b11110110110001110001101100000000;
   assign mem[72703:72672] = 32'b00001100010011111010100011110000;
   assign mem[72735:72704] = 32'b11101011000000000010110011000000;
   assign mem[72767:72736] = 32'b00000001101111111111010100000110;
   assign mem[72799:72768] = 32'b00001100110111010011100111010000;
   assign mem[72831:72800] = 32'b11111110100000011011010011101000;
   assign mem[72863:72832] = 32'b00000110111000011001111001111000;
   assign mem[72895:72864] = 32'b11100100111001010011000001000000;
   assign mem[72927:72896] = 32'b00000010111001011010110110000000;
   assign mem[72959:72928] = 32'b11110001011101111101111101110000;
   assign mem[72991:72960] = 32'b11111100111101110011011111100100;
   assign mem[73023:72992] = 32'b00000000101000010000000001101100;
   assign mem[73055:73024] = 32'b11111111011011111111100100100010;
   assign mem[73087:73056] = 32'b00000010100000000100100110101000;
   assign mem[73119:73088] = 32'b11111010111000111111000000110000;
   assign mem[73151:73120] = 32'b11111110000010111101000100100010;
   assign mem[73183:73152] = 32'b11111010100101110010101101111000;
   assign mem[73215:73184] = 32'b11111110001110001010010101110010;
   assign mem[73247:73216] = 32'b00000001010001100001110111111100;
   assign mem[73279:73248] = 32'b00000100001001111111101010101000;
   assign mem[73311:73280] = 32'b11111111000111110110010001100010;
   assign mem[73343:73312] = 32'b11111110001010110000100111010010;
   assign mem[73375:73344] = 32'b00000010100100011101100100111100;
   assign mem[73407:73376] = 32'b00000000110100011110011101011111;
   assign mem[73439:73408] = 32'b11111100001111011000001101001000;
   assign mem[73471:73440] = 32'b11111100110000000111110001101100;
   assign mem[73503:73472] = 32'b11111001101111110101001101010000;
   assign mem[73535:73504] = 32'b00000110001001110001100001011000;
   assign mem[73567:73536] = 32'b00000010101001011101111011010100;
   assign mem[73599:73568] = 32'b00000101010001101010101100110000;
   assign mem[73631:73600] = 32'b11111100011000000101111101000100;
   assign mem[73663:73632] = 32'b00000001100000000101000100101000;
   assign mem[73695:73664] = 32'b11111001011111001000101010001000;
   assign mem[73727:73696] = 32'b11111110000101111110100101011100;
   assign mem[73759:73728] = 32'b00000001010000111111011011001100;
   assign mem[73791:73760] = 32'b00000110101111111111100010111000;
   assign mem[73823:73792] = 32'b11111110111111000010101111101000;
   assign mem[73855:73824] = 32'b00000001001001111100000111111000;
   assign mem[73887:73856] = 32'b00000010001011000101001001010000;
   assign mem[73919:73888] = 32'b11111000011001111010101010101000;
   assign mem[73951:73920] = 32'b11111100111101001101100101100100;
   assign mem[73983:73952] = 32'b00000010011011111000010001100100;
   assign mem[74015:73984] = 32'b11101111001010001101110101100000;
   assign mem[74047:74016] = 32'b11111001101100001100111001111000;
   assign mem[74079:74048] = 32'b00000100100010111001111100110000;
   assign mem[74111:74080] = 32'b00000100111011010101010110110000;
   assign mem[74143:74112] = 32'b11111101011001101001110001010100;
   assign mem[74175:74144] = 32'b00000000011010011101001011000110;
   assign mem[74207:74176] = 32'b11111001000011010011111010000000;
   assign mem[74239:74208] = 32'b00000011100000011101010110001000;
   assign mem[74271:74240] = 32'b00000000000000101000110111000100;
   assign mem[74303:74272] = 32'b11111010110011011010000111001000;
   assign mem[74335:74304] = 32'b00001000010101010011011101000000;
   assign mem[74367:74336] = 32'b00000000111010100000110001010010;
   assign mem[74399:74368] = 32'b11111010100100000011000100010000;
   assign mem[74431:74400] = 32'b11111011010100100011101110100000;
   assign mem[74463:74432] = 32'b11111111100100110011101110011101;
   assign mem[74495:74464] = 32'b11111110110001011000001111000100;
   assign mem[74527:74496] = 32'b11110011100011001110011100110000;
   assign mem[74559:74528] = 32'b00000100110101001100100111100000;
   assign mem[74591:74560] = 32'b11111100000111010101100011011000;
   assign mem[74623:74592] = 32'b00000011010000010110001100100100;
   assign mem[74655:74624] = 32'b11110111100011010001010110000000;
   assign mem[74687:74656] = 32'b11111100101011011110000111001000;
   assign mem[74719:74688] = 32'b11101110010011011001000010100000;
   assign mem[74751:74720] = 32'b00001001000101011110111100110000;
   assign mem[74783:74752] = 32'b00000001001110010100000101100010;
   assign mem[74815:74784] = 32'b11110111100010111101100111100000;
   assign mem[74847:74816] = 32'b00000001100100011010000100100100;
   assign mem[74879:74848] = 32'b00000100110011000101101101000000;
   assign mem[74911:74880] = 32'b11111111000110111100111010011111;
   assign mem[74943:74912] = 32'b11111111111010100011001111000010;
   assign mem[74975:74944] = 32'b11111100010101011100011000010000;
   assign mem[75007:74976] = 32'b00000100100110101111000010000000;
   assign mem[75039:75008] = 32'b11110100011011111000001101010000;
   assign mem[75071:75040] = 32'b00000010111100011001000001011100;
   assign mem[75103:75072] = 32'b11111111001110011001010110000010;
   assign mem[75135:75104] = 32'b00001001001101101001100010110000;
   assign mem[75167:75136] = 32'b11110100100000000101110010000000;
   assign mem[75199:75168] = 32'b11101111101011010100100101000000;
   assign mem[75231:75200] = 32'b11111010101111010000011100010000;
   assign mem[75263:75232] = 32'b00000010100010111110010110010100;
   assign mem[75295:75264] = 32'b00000011101111001111110000100100;
   assign mem[75327:75296] = 32'b00000110011010100100100011100000;
   assign mem[75359:75328] = 32'b00001000001101001001101010000000;
   assign mem[75391:75360] = 32'b11110110111011011001000001000000;
   assign mem[75423:75392] = 32'b11111011111100110001111110101000;
   assign mem[75455:75424] = 32'b00000010100011010001011100100100;
   assign mem[75487:75456] = 32'b00000000000111001011000101111000;
   assign mem[75519:75488] = 32'b11111000100000001000001111111000;
   assign mem[75551:75520] = 32'b11111011000001010101110011101000;
   assign mem[75583:75552] = 32'b00000010001000111010001100100100;
   assign mem[75615:75584] = 32'b11111100000010101001000010000100;
   assign mem[75647:75616] = 32'b00000010001100100001000111110000;
   assign mem[75679:75648] = 32'b00000101101010010110100000100000;
   assign mem[75711:75680] = 32'b00000001001010110011000000111110;
   assign mem[75743:75712] = 32'b11110110111101011010111100110000;
   assign mem[75775:75744] = 32'b00000010000100100101101101110100;
   assign mem[75807:75776] = 32'b00000010000110010001000001010100;
   assign mem[75839:75808] = 32'b11111110011110110111110011011110;
   assign mem[75871:75840] = 32'b00000001100100001001010010011010;
   assign mem[75903:75872] = 32'b11111001011111100011101111111000;
   assign mem[75935:75904] = 32'b00000010110101011111111110111100;
   assign mem[75967:75936] = 32'b00000101010110101001101000010000;
   assign mem[75999:75968] = 32'b11111000111101110010011011100000;
   assign mem[76031:76000] = 32'b11110110011001000000001010000000;
   assign mem[76063:76032] = 32'b11111101010000101010111000100100;
   assign mem[76095:76064] = 32'b00000010100111100011011000011100;
   assign mem[76127:76096] = 32'b00000011100010000100000111000100;
   assign mem[76159:76128] = 32'b00000100011011111000101001001000;
   assign mem[76191:76160] = 32'b11111110010010001100010100010010;
   assign mem[76223:76192] = 32'b00000100101100010001111111011000;
   assign mem[76255:76224] = 32'b00000101011010001000100010101000;
   assign mem[76287:76256] = 32'b00000010000110111111010110101100;
   assign mem[76319:76288] = 32'b00000000010011101100001011100001;
   assign mem[76351:76320] = 32'b00000001110011110100001000011100;
   assign mem[76383:76352] = 32'b11110101111001010001101000010000;
   assign mem[76415:76384] = 32'b11110010011100101001010111000000;
   assign mem[76447:76416] = 32'b11111000001000001110010000000000;
   assign mem[76479:76448] = 32'b11111011010010001010101010000000;
   assign mem[76511:76480] = 32'b11111110110010011001101101100000;
   assign mem[76543:76512] = 32'b00000010100110011001100111011000;
   assign mem[76575:76544] = 32'b11111100111010001100100011111100;
   assign mem[76607:76576] = 32'b11111100101011000000010000000100;
   assign mem[76639:76608] = 32'b00000011000010011100001000110100;
   assign mem[76671:76640] = 32'b11111101001011001000011110011100;
   assign mem[76703:76672] = 32'b00000001101100101010110000110110;
   assign mem[76735:76704] = 32'b00000010011101111111100100001100;
   assign mem[76767:76736] = 32'b11111111110001001010011000010011;
   assign mem[76799:76768] = 32'b11111100001111100101110110000100;
   assign mem[76831:76800] = 32'b00000100001011101000010111100000;
   assign mem[76863:76832] = 32'b11110011110100110110011010010000;
   assign mem[76895:76864] = 32'b11111110010010010011001000101010;
   assign mem[76927:76896] = 32'b00000000101101111111010011011001;
   assign mem[76959:76928] = 32'b11110011111101011111001101000000;
   assign mem[76991:76960] = 32'b00000111001001001010010010100000;
   assign mem[77023:76992] = 32'b00000011100100101001001000111000;
   assign mem[77055:77024] = 32'b11111000101100001111100000011000;
   assign mem[77087:77056] = 32'b00000001111000100011000010100000;
   assign mem[77119:77088] = 32'b11111001110100000010111111100000;
   assign mem[77151:77120] = 32'b11111111101100100100111000011010;
   assign mem[77183:77152] = 32'b00000100010011001011001101111000;
   assign mem[77215:77184] = 32'b11111011111001111001101011111000;
   assign mem[77247:77216] = 32'b11110110011100011100111000110000;
   assign mem[77279:77248] = 32'b00000011101001000011111110100100;
   assign mem[77311:77280] = 32'b00000101010011010011101001001000;
   assign mem[77343:77312] = 32'b00000001001101011000001001001000;
   assign mem[77375:77344] = 32'b11111011010000111111010010000000;
   assign mem[77407:77376] = 32'b11111011010110011111000110000000;
   assign mem[77439:77408] = 32'b00000010101010110001111110110000;
   assign mem[77471:77440] = 32'b11111110100010000111101011101100;
   assign mem[77503:77472] = 32'b00000010110001011110110101111100;
   assign mem[77535:77504] = 32'b00000000001001101100101011000011;
   assign mem[77567:77536] = 32'b11111110100001010011000010000100;
   assign mem[77599:77568] = 32'b00000100011110100001000101101000;
   assign mem[77631:77600] = 32'b00000001010001110100100100000100;
   assign mem[77663:77632] = 32'b00000100100010111101000101110000;
   assign mem[77695:77664] = 32'b11111001101001001100100100110000;
   assign mem[77727:77696] = 32'b11111111110001011000111101000100;
   assign mem[77759:77728] = 32'b11111100111111101100110111000000;
   assign mem[77791:77760] = 32'b00000000000111001110101110101010;
   assign mem[77823:77792] = 32'b00001010110110111110111001010000;
   assign mem[77855:77824] = 32'b11110110111001010100110111010000;
   assign mem[77887:77856] = 32'b11111100101100100111010011011100;
   assign mem[77919:77888] = 32'b00001000100110101001001000110000;
   assign mem[77951:77920] = 32'b11110111100111011111110000000000;
   assign mem[77983:77952] = 32'b00001101011001100000100010000000;
   assign mem[78015:77984] = 32'b11111110000011001011100011010110;
   assign mem[78047:78016] = 32'b00000011110010010100100111001100;
   assign mem[78079:78048] = 32'b11110101111001000100101110010000;
   assign mem[78111:78080] = 32'b00000011101111110111101000000000;
   assign mem[78143:78112] = 32'b11111011111011110010010010000000;
   assign mem[78175:78144] = 32'b11111110000011100011101101100000;
   assign mem[78207:78176] = 32'b00000101010111011111011010000000;
   assign mem[78239:78208] = 32'b11100110011001010010001010100000;
   assign mem[78271:78240] = 32'b00000100100001111111001100000000;
   assign mem[78303:78272] = 32'b00000001111000101011001110101010;
   assign mem[78335:78304] = 32'b11111011111100100011000100111000;
   assign mem[78367:78336] = 32'b00000001010001100100001000011100;
   assign mem[78399:78368] = 32'b00000010111000011101001010111000;
   assign mem[78431:78400] = 32'b00000001001000111001011001001000;
   assign mem[78463:78432] = 32'b11101111110011110100111011000000;
   assign mem[78495:78464] = 32'b11111111111010011000011101110100;
   assign mem[78527:78496] = 32'b00000000010111100010111010100110;
   assign mem[78559:78528] = 32'b11110001000011110110101100100000;
   assign mem[78591:78560] = 32'b00000100010100001010100111000000;
   assign mem[78623:78592] = 32'b11111101001101101001110110101100;
   assign mem[78655:78624] = 32'b00000101001001100110001011010000;
   assign mem[78687:78656] = 32'b00000000010001011000101111010000;
   assign mem[78719:78688] = 32'b00000111011111011000011000001000;
   assign mem[78751:78720] = 32'b11111111001101000000100111010011;
   assign mem[78783:78752] = 32'b11111111101001101010101100000011;
   assign mem[78815:78784] = 32'b11111101011000000110111000000100;
   assign mem[78847:78816] = 32'b11111100011010100000101010101100;
   assign mem[78879:78848] = 32'b11110001100001100000101100100000;
   assign mem[78911:78880] = 32'b00000111010101100010101000001000;
   assign mem[78943:78912] = 32'b00000110100111101001000011111000;
   assign mem[78975:78944] = 32'b11101101010010110011010110100000;
   assign mem[79007:78976] = 32'b11111101011000110100111010110000;
   assign mem[79039:79008] = 32'b00000100001001110100110001100000;
   assign mem[79071:79040] = 32'b11110101100010110001100101010000;
   assign mem[79103:79072] = 32'b00000100010000111000111000010000;
   assign mem[79135:79104] = 32'b11110001110011100011000101010000;
   assign mem[79167:79136] = 32'b00000001100100111010010010011010;
   assign mem[79199:79168] = 32'b00010000001101111000011101100000;
   assign mem[79231:79200] = 32'b00000010100111010100111010000000;
   assign mem[79263:79232] = 32'b00000101101010010111101001001000;
   assign mem[79295:79264] = 32'b11110101100111000111101110000000;
   assign mem[79327:79296] = 32'b00000001000001010101110100101110;
   assign mem[79359:79328] = 32'b11101110100010101010001001100000;
   assign mem[79391:79360] = 32'b11111111110010110001111101110011;
   assign mem[79423:79392] = 32'b00000010011101001101101011000100;
   assign mem[79455:79424] = 32'b00000001110101101100101001011110;
   assign mem[79487:79456] = 32'b00001011110101100100000000010000;
   assign mem[79519:79488] = 32'b11111110001100001100011111001110;
   assign mem[79551:79520] = 32'b11110110110101100010101111110000;
   assign mem[79583:79552] = 32'b11111101001111000110110100110000;
   assign mem[79615:79584] = 32'b00000010111110011100111001000000;
   assign mem[79647:79616] = 32'b11111110000011101101110111001110;
   assign mem[79679:79648] = 32'b11110100011011101001111010010000;
   assign mem[79711:79680] = 32'b00000011000100110110110011110100;
   assign mem[79743:79712] = 32'b11110011011100011110010000100000;
   assign mem[79775:79744] = 32'b00000101001101011011000001110000;
   assign mem[79807:79776] = 32'b00001100001010010001001110110000;
   assign mem[79839:79808] = 32'b11111101111101100111001010100100;
   assign mem[79871:79840] = 32'b11111101101111011111111000110000;
   assign mem[79903:79872] = 32'b11111011010110101101111111011000;
   assign mem[79935:79904] = 32'b11111100011001110000100111100100;
   assign mem[79967:79936] = 32'b11111100111000011111101011010100;
   assign mem[79999:79968] = 32'b11111010111110110011001011011000;
   assign mem[80031:80000] = 32'b00000000000111010101010111100011;
   assign mem[80063:80032] = 32'b00000001100110000100001101110000;
   assign mem[80095:80064] = 32'b11111100111011000111011011111000;
   assign mem[80127:80096] = 32'b00000000001100000101111001100111;
   assign mem[80159:80128] = 32'b11111101010000000010110111101000;
   assign mem[80191:80160] = 32'b11111111011011001011100111111100;
   assign mem[80223:80192] = 32'b11111001001000111111011100100000;
   assign mem[80255:80224] = 32'b11111111001100110111110011010001;
   assign mem[80287:80256] = 32'b11111111011110100011101011011111;
   assign mem[80319:80288] = 32'b11111111111010010110001011100010;
   assign mem[80351:80320] = 32'b00000011010001011101101100100000;
   assign mem[80383:80352] = 32'b11111111011100000100000001111111;
   assign mem[80415:80384] = 32'b00000010001001101110010001110100;
   assign mem[80447:80416] = 32'b11111111011000100011011000011110;
   assign mem[80479:80448] = 32'b11111111010000010100100111101111;
   assign mem[80511:80480] = 32'b11111110111111010101101010101100;
   assign mem[80543:80512] = 32'b11110110100101111011011001100000;
   assign mem[80575:80544] = 32'b11111111001011010110111101111101;
   assign mem[80607:80576] = 32'b00000001001100101011100011011110;
   assign mem[80639:80608] = 32'b00000010010011110111100000001000;
   assign mem[80671:80640] = 32'b00000000110101111011101000110100;
   assign mem[80703:80672] = 32'b00000100100010100101111010001000;
   assign mem[80735:80704] = 32'b00000000010111100010001010010110;
   assign mem[80767:80736] = 32'b11111100110001001100110110100100;
   assign mem[80799:80768] = 32'b00000101000010111000001101001000;
   assign mem[80831:80800] = 32'b00000000001010001000001010010111;
   assign mem[80863:80832] = 32'b11111111011100001110100101001010;
   assign mem[80895:80864] = 32'b11111111100110001100110000101100;
   assign mem[80927:80896] = 32'b00000001010011011011101001100000;
   assign mem[80959:80928] = 32'b00000010011110100011000010011100;
   assign mem[80991:80960] = 32'b00000100010101000101101011010000;
   assign mem[81023:80992] = 32'b00000101010010101000100111010000;
   assign mem[81055:81024] = 32'b11111010100100010011000100110000;
   assign mem[81087:81056] = 32'b11110110000001010101100011110000;
   assign mem[81119:81088] = 32'b00000100010110110000011000111000;
   assign mem[81151:81120] = 32'b11111101011001111100110101001000;
   assign mem[81183:81152] = 32'b00000001001001101101010100010110;
   assign mem[81215:81184] = 32'b00000010110111000101000001111100;
   assign mem[81247:81216] = 32'b11111101000111111010110110110100;
   assign mem[81279:81248] = 32'b00000001000001000110000010110110;
   assign mem[81311:81280] = 32'b11111011111100011100100100101000;
   assign mem[81343:81312] = 32'b00000011011111000101001111110100;
   assign mem[81375:81344] = 32'b00000011010000001110011011100100;
   assign mem[81407:81376] = 32'b11110110001011000001110001110000;
   assign mem[81439:81408] = 32'b00001110101100101100001101010000;
   assign mem[81471:81440] = 32'b11111111000101001101111101110101;
   assign mem[81503:81472] = 32'b00000011001110001111101001110100;
   assign mem[81535:81504] = 32'b11101110110010000111111100000000;
   assign mem[81567:81536] = 32'b00000000010110101111110101111001;
   assign mem[81599:81568] = 32'b11101010001001100100010110100000;
   assign mem[81631:81600] = 32'b11111101111000001111011010100100;
   assign mem[81663:81632] = 32'b00001001011001000001110001000000;
   assign mem[81695:81664] = 32'b11111000010101011001110100110000;
   assign mem[81727:81696] = 32'b00000000011001111010111101001111;
   assign mem[81759:81728] = 32'b00001001110001000111001000100000;
   assign mem[81791:81760] = 32'b00000101010101111100111010011000;
   assign mem[81823:81792] = 32'b00000000101000000110100001010011;
   assign mem[81855:81824] = 32'b11111111000000000100111101010001;
   assign mem[81887:81856] = 32'b11111111001001100000111101001011;
   assign mem[81919:81888] = 32'b11110100011101001110101011000000;
   assign mem[81951:81920] = 32'b00000101000110100000001100111000;
   assign mem[81983:81952] = 32'b11111001101110110100011000111000;
   assign mem[82015:81984] = 32'b11110101011101110110101011110000;
   assign mem[82047:82016] = 32'b11111101000101111110111110011000;
   assign mem[82079:82048] = 32'b11111111010001101011011011011101;
   assign mem[82111:82080] = 32'b11111110111010010010110110011110;
   assign mem[82143:82112] = 32'b11111101111110001001100011011100;
   assign mem[82175:82144] = 32'b00000100101011111011100000010000;
   assign mem[82207:82176] = 32'b00000101101010000110000111101000;
   assign mem[82239:82208] = 32'b00000011011000011010101110100100;
   assign mem[82271:82240] = 32'b11111110110110011010001000001000;
   assign mem[82303:82272] = 32'b00000000101110101011110010010011;
   assign mem[82335:82304] = 32'b11111110101000011110110110110100;
   assign mem[82367:82336] = 32'b00000000011000001100111001010011;
   assign mem[82399:82368] = 32'b00000000000010010010111101011100;
   assign mem[82431:82400] = 32'b11111000001100010111000001011000;
   assign mem[82463:82432] = 32'b11111001100111110111111111111000;
   assign mem[82495:82464] = 32'b11111110011010011001000100010000;
   assign mem[82527:82496] = 32'b00000000101001011110100011101010;
   assign mem[82559:82528] = 32'b00000010000011111010101001110000;
   assign mem[82591:82560] = 32'b00000101100111000110001100100000;
   assign mem[82623:82592] = 32'b11110100101011011011010101000000;
   assign mem[82655:82624] = 32'b00000011000000111001111111101000;
   assign mem[82687:82656] = 32'b00000111110111010100111100011000;
   assign mem[82719:82688] = 32'b11111001110001000110001001001000;
   assign mem[82751:82720] = 32'b11110000101101111110000001110000;
   assign mem[82783:82752] = 32'b00000110011011110000011100100000;
   assign mem[82815:82784] = 32'b00000010111100111101011010010100;
   assign mem[82847:82816] = 32'b00000001111110011010010000011110;
   assign mem[82879:82848] = 32'b00000100001010010001000101100000;
   assign mem[82911:82880] = 32'b11111100101101101100110101101000;
   assign mem[82943:82912] = 32'b11110101001011000010010111010000;
   assign mem[82975:82944] = 32'b11111000010001000111110000001000;
   assign mem[83007:82976] = 32'b11110010100011000001011000010000;
   assign mem[83039:83008] = 32'b11111101110101000111110110011000;
   assign mem[83071:83040] = 32'b00000010101001101010010101010000;
   assign mem[83103:83072] = 32'b11111110011011101110001101100010;
   assign mem[83135:83104] = 32'b11110001111001111100111110010000;
   assign mem[83167:83136] = 32'b00000011000010110001110100010000;
   assign mem[83199:83168] = 32'b11110101011010011011101100000000;
   assign mem[83231:83200] = 32'b11111010011000010010111110000000;
   assign mem[83263:83232] = 32'b00000000010001110110010010000000;
   assign mem[83295:83264] = 32'b11110110001000000001010001010000;
   assign mem[83327:83296] = 32'b11101100010010000011011111000000;
   assign mem[83359:83328] = 32'b11111100101111000001111011111000;
   assign mem[83391:83360] = 32'b00000101001111110000110011011000;
   assign mem[83423:83392] = 32'b00001001101010100001101110010000;
   assign mem[83455:83424] = 32'b11111100011011011010000001001100;
   assign mem[83487:83456] = 32'b11111111011000010001000100110010;
   assign mem[83519:83488] = 32'b11111011001110001111111010101000;
   assign mem[83551:83520] = 32'b00000111111100000101100101001000;
   assign mem[83583:83552] = 32'b00000111111110111010100011111000;
   assign mem[83615:83584] = 32'b11111001011011100001010101111000;
   assign mem[83647:83616] = 32'b11110110111001011000001011110000;
   assign mem[83679:83648] = 32'b00000111110001010111111110000000;
   assign mem[83711:83680] = 32'b00000010000110000100000101011100;
   assign mem[83743:83712] = 32'b00000010111010010101111010101000;
   assign mem[83775:83744] = 32'b11111111110011011000001001010000;
   assign mem[83807:83776] = 32'b11111101101000000000000000010100;
   assign mem[83839:83808] = 32'b11110110110010001110110001010000;
   assign mem[83871:83840] = 32'b11110011110111111000001001010000;
   assign mem[83903:83872] = 32'b11111111100011100100111111111101;
   assign mem[83935:83904] = 32'b11111101011100001110010011000000;
   assign mem[83967:83936] = 32'b00000011010111000101000001001100;
   assign mem[83999:83968] = 32'b11111010100111100100010000100000;
   assign mem[84031:84000] = 32'b00000001010101001111001011110100;
   assign mem[84063:84032] = 32'b00000011011011100100111100011000;
   assign mem[84095:84064] = 32'b00000010011011111001101100100100;
   assign mem[84127:84096] = 32'b00000000111001111110111111111010;
   assign mem[84159:84128] = 32'b11111000010100000000100010111000;
   assign mem[84191:84160] = 32'b11110110111101010011110000110000;
   assign mem[84223:84192] = 32'b00001001111000001010011011100000;
   assign mem[84255:84224] = 32'b11101100011010101010011011100000;
   assign mem[84287:84256] = 32'b11111011111011101111110110000000;
   assign mem[84319:84288] = 32'b00000001001101101010100100001010;
   assign mem[84351:84320] = 32'b00001001010011001001110100010000;
   assign mem[84383:84352] = 32'b00000100010010100101010001110000;
   assign mem[84415:84384] = 32'b00000011001100101101100101001100;
   assign mem[84447:84416] = 32'b11111110011011110101111001000010;
   assign mem[84479:84448] = 32'b00000010000000001110011111100100;
   assign mem[84511:84480] = 32'b11111110101010111111101110111010;
   assign mem[84543:84512] = 32'b00000000010000011001100101010100;
   assign mem[84575:84544] = 32'b11111011111010001110001010100000;
   assign mem[84607:84576] = 32'b11111101111110001001011000010000;
   assign mem[84639:84608] = 32'b11111111111011110011001000111000;
   assign mem[84671:84640] = 32'b11111111001010101010110001101010;
   assign mem[84703:84672] = 32'b11111110010011000101001110001000;
   assign mem[84735:84704] = 32'b00000011001100001101111110000000;
   assign mem[84767:84736] = 32'b00000010011000000100110111010000;
   assign mem[84799:84768] = 32'b00000001100110011011111000010000;
   assign mem[84831:84800] = 32'b11101000110111101011011010000000;
   assign mem[84863:84832] = 32'b00001010101110111111010001110000;
   assign mem[84895:84864] = 32'b11110001101101110111100111000000;
   assign mem[84927:84896] = 32'b11111001110110010011010111010000;
   assign mem[84959:84928] = 32'b00000101110111110100101010010000;
   assign mem[84991:84960] = 32'b00001011011100111001111001000000;
   assign mem[85023:84992] = 32'b00010001000111111000101110000000;
   assign mem[85055:85024] = 32'b11111111001001101010111000000000;
   assign mem[85087:85056] = 32'b11111011110001001110011101101000;
   assign mem[85119:85088] = 32'b11110010111100001101100100110000;
   assign mem[85151:85120] = 32'b11111101100010110111011010100100;
   assign mem[85183:85152] = 32'b11111101001100000111010000010000;
   assign mem[85215:85184] = 32'b11111110001010111101000101111110;
   assign mem[85247:85216] = 32'b00000000000101101010111001010110;
   assign mem[85279:85248] = 32'b00000011010000111001111111001100;
   assign mem[85311:85280] = 32'b00000100111100100100100001010000;
   assign mem[85343:85312] = 32'b00000010010011111001011000011100;
   assign mem[85375:85344] = 32'b00000001011000110110101110000110;
   assign mem[85407:85376] = 32'b11111111111111101111011000100111;
   assign mem[85439:85408] = 32'b00000010001010011101111010111100;
   assign mem[85471:85440] = 32'b11111111000101110000000101000000;
   assign mem[85503:85472] = 32'b11111011111100001011011000100000;
   assign mem[85535:85504] = 32'b00000010110011000110011111001100;
   assign mem[85567:85536] = 32'b00000001011000110000001110010110;
   assign mem[85599:85568] = 32'b11110110101111101011100001010000;
   assign mem[85631:85600] = 32'b11111000011100001100000111011000;
   assign mem[85663:85632] = 32'b00001001000100100110010100010000;
   assign mem[85695:85664] = 32'b11111010001110010100100001000000;
   assign mem[85727:85696] = 32'b00000101011001010100011101100000;
   assign mem[85759:85728] = 32'b11111100010100100110001011101000;
   assign mem[85791:85760] = 32'b11111101100000011010011001001000;
   assign mem[85823:85792] = 32'b11111111010011101110000010011001;
   assign mem[85855:85824] = 32'b11111011001011010011100000001000;
   assign mem[85887:85856] = 32'b11111111000011100010000101111000;
   assign mem[85919:85888] = 32'b11111001100000000101000101101000;
   assign mem[85951:85920] = 32'b00000100110110000000011111110000;
   assign mem[85983:85952] = 32'b11111001111000100110001000101000;
   assign mem[86015:85984] = 32'b00000110001011111011010011000000;
   assign mem[86047:86016] = 32'b00000100011001110010100000001000;
   assign mem[86079:86048] = 32'b00000010001111100101111100110100;
   assign mem[86111:86080] = 32'b00000010011011000001110001001100;
   assign mem[86143:86112] = 32'b11111011100001001101110011010000;
   assign mem[86175:86144] = 32'b11111101100111101101110011110000;
   assign mem[86207:86176] = 32'b11111100101010110111110001100000;
   assign mem[86239:86208] = 32'b11111110001000010110010001101000;
   assign mem[86271:86240] = 32'b00000001001011110010010111000010;
   assign mem[86303:86272] = 32'b11111111011010111100101000000110;
   assign mem[86335:86304] = 32'b00000000110010011010011101001001;
   assign mem[86367:86336] = 32'b00000001100111001001111110000110;
   assign mem[86399:86368] = 32'b00000000001000110111001110111110;
   assign mem[86431:86400] = 32'b00001000000100101101001011110000;
   assign mem[86463:86432] = 32'b11111011110011000011110001111000;
   assign mem[86495:86464] = 32'b00000010010010010011001000110000;
   assign mem[86527:86496] = 32'b00000010110000100110010001001100;
   assign mem[86559:86528] = 32'b11110110100111001010001111000000;
   assign mem[86591:86560] = 32'b00000100100010000110101001000000;
   assign mem[86623:86592] = 32'b11111100001001100010111110000100;
   assign mem[86655:86624] = 32'b00001011000010001011000110110000;
   assign mem[86687:86656] = 32'b11111111010111000100100001111100;
   assign mem[86719:86688] = 32'b11111100111000111001110010101000;
   assign mem[86751:86720] = 32'b11111100011001110000110011000100;
   assign mem[86783:86752] = 32'b00001010101100001011101111000000;
   assign mem[86815:86784] = 32'b11101010100110110011111110100000;
   assign mem[86847:86816] = 32'b11100000011111101011010011100000;
   assign mem[86879:86848] = 32'b00001010011010001100000100110000;
   assign mem[86911:86880] = 32'b00001001100001111010010000010000;
   assign mem[86943:86912] = 32'b00000011000100110001000000001100;
   assign mem[86975:86944] = 32'b11110101111011110101100111010000;
   assign mem[87007:86976] = 32'b00001001000101101101001100110000;
   assign mem[87039:87008] = 32'b11101000000101111010110100000000;
   assign mem[87071:87040] = 32'b11111110010111111011000110011010;
   assign mem[87103:87072] = 32'b11111101110000010100110100000100;
   assign mem[87135:87104] = 32'b11101110101100100111111110000000;
   assign mem[87167:87136] = 32'b11101111011101011101000111100000;
   assign mem[87199:87168] = 32'b11111011010011010100110001000000;
   assign mem[87231:87200] = 32'b00001010000010000111100110100000;
   assign mem[87263:87232] = 32'b00000000011111111110001010111000;
   assign mem[87295:87264] = 32'b11110010100000001100101100010000;
   assign mem[87327:87296] = 32'b00000110110000111111001100101000;
   assign mem[87359:87328] = 32'b11111001011100001100111000110000;
   assign mem[87391:87360] = 32'b00000010100100001110011011001000;
   assign mem[87423:87392] = 32'b11101111011000100111111010100000;
   assign mem[87455:87424] = 32'b00000111000010110101111111010000;
   assign mem[87487:87456] = 32'b00000110111010101011011011110000;
   assign mem[87519:87488] = 32'b11110000101011111110100001110000;
   assign mem[87551:87520] = 32'b11111000111100111111010000010000;
   assign mem[87583:87552] = 32'b11111111101010101011011011101110;
   assign mem[87615:87584] = 32'b00000000001110011101010000100111;
   assign mem[87647:87616] = 32'b00000000110101000110110110100110;
   assign mem[87679:87648] = 32'b00000011111101011101000110010000;
   assign mem[87711:87680] = 32'b00000101111111101010111010011000;
   assign mem[87743:87712] = 32'b11111110100111010101000101000110;
   assign mem[87775:87744] = 32'b11111111000111110011100110101111;
   assign mem[87807:87776] = 32'b11111111011010111110001101110101;
   assign mem[87839:87808] = 32'b11111111011001000111100110111101;
   assign mem[87871:87840] = 32'b11111010111101000111000111110000;
   assign mem[87903:87872] = 32'b11110111101010100000011011010000;
   assign mem[87935:87904] = 32'b11111111010010011100011010110110;
   assign mem[87967:87936] = 32'b00000011111011101010011101010000;
   assign mem[87999:87968] = 32'b00000010001100111010000110100100;
   assign mem[88031:88000] = 32'b00000001101011110100000111000000;
   assign mem[88063:88032] = 32'b11111110000011011111010111000110;
   assign mem[88095:88064] = 32'b11110011110011100101100010110000;
   assign mem[88127:88096] = 32'b11111110110000000111101011101100;
   assign mem[88159:88128] = 32'b00000001101011000111001110100110;
   assign mem[88191:88160] = 32'b00000100110101110001001100011000;
   assign mem[88223:88192] = 32'b11111101000100001110001000001100;
   assign mem[88255:88224] = 32'b00000010011110111001010010110100;
   assign mem[88287:88256] = 32'b11111110100010000110110101111110;
   assign mem[88319:88288] = 32'b00000100010100000000101010011000;
   assign mem[88351:88320] = 32'b11111011001110111111111100111000;
   assign mem[88383:88352] = 32'b00000010100011110010001111000000;
   assign mem[88415:88384] = 32'b11111000011010101110000100110000;
   assign mem[88447:88416] = 32'b11110101010101010010100111000000;
   assign mem[88479:88448] = 32'b00000011101101111011111101101100;
   assign mem[88511:88480] = 32'b00000000101000101000111111001010;
   assign mem[88543:88512] = 32'b11111101001101000010101000110000;
   assign mem[88575:88544] = 32'b11111110110101101011010110000010;
   assign mem[88607:88576] = 32'b00000100101000111110000101100000;
   assign mem[88639:88608] = 32'b11111001111000100100001110111000;
   assign mem[88671:88640] = 32'b00000001101101010111101111110000;
   assign mem[88703:88672] = 32'b11111100101010000000000011100000;
   assign mem[88735:88704] = 32'b11111100001100111101111101000000;
   assign mem[88767:88736] = 32'b11111110100010001001101101011110;
   assign mem[88799:88768] = 32'b00000101111011110010111011110000;
   assign mem[88831:88800] = 32'b00001000011101000111100101110000;
   assign mem[88863:88832] = 32'b11111100110111111100100110111100;
   assign mem[88895:88864] = 32'b00000010100010101100111100001000;
   assign mem[88927:88896] = 32'b11111111001000110000111111110100;
   assign mem[88959:88928] = 32'b11111111110011010011100010110101;
   assign mem[88991:88960] = 32'b11111110101000111110001111111000;
   assign mem[89023:88992] = 32'b00000110100110111010111000001000;
   assign mem[89055:89024] = 32'b11101110000011011001001101000000;
   assign mem[89087:89056] = 32'b00000010011011111000010001111000;
   assign mem[89119:89088] = 32'b00000101000011111100000101100000;
   assign mem[89151:89120] = 32'b00000010000001010010010000100000;
   assign mem[89183:89152] = 32'b00000110100001011101110000111000;
   assign mem[89215:89184] = 32'b00000101000010001011110100111000;
   assign mem[89247:89216] = 32'b00000010011011001101111100011100;
   assign mem[89279:89248] = 32'b11110101001000101000101100010000;
   assign mem[89311:89280] = 32'b00000011100111111111100111000000;
   assign mem[89343:89312] = 32'b11110111111101100101000111110000;
   assign mem[89375:89344] = 32'b00000011000000001000110101101100;
   assign mem[89407:89376] = 32'b00000001111010001001001011000110;
   assign mem[89439:89408] = 32'b00000010111001010111111101001100;
   assign mem[89471:89440] = 32'b11110000010000001010011111010000;
   assign mem[89503:89472] = 32'b00000001011110011100111000100010;
   assign mem[89535:89504] = 32'b11111101111000110110001011101100;
   assign mem[89567:89536] = 32'b00000000110111011111000100111111;
   assign mem[89599:89568] = 32'b00000000010100011011001111001011;
   assign mem[89631:89600] = 32'b00000100001011110000001001011000;
   assign mem[89663:89632] = 32'b00000110110001110010001011011000;
   assign mem[89695:89664] = 32'b11111101100110101010100000100100;
   assign mem[89727:89696] = 32'b00000000001110010001001011001101;
   assign mem[89759:89728] = 32'b00000001001010011001010001110100;
   assign mem[89791:89760] = 32'b11101110011110110110100110000000;
   assign mem[89823:89792] = 32'b00000101110111110010111010110000;
   assign mem[89855:89824] = 32'b11111010111001000001100000101000;
   assign mem[89887:89856] = 32'b00000100111110100100011000110000;
   assign mem[89919:89888] = 32'b11110110101010110110111101100000;
   assign mem[89951:89920] = 32'b11111010110000000100000101111000;
   assign mem[89983:89952] = 32'b00000110101110001011100110101000;
   assign mem[90015:89984] = 32'b00000100010000101101010101001000;
   assign mem[90047:90016] = 32'b00000011110100100001010100010100;
   assign mem[90079:90048] = 32'b11111100101101000100101100100100;
   assign mem[90111:90080] = 32'b11111101100111011011110101010100;
   assign mem[90143:90112] = 32'b11111110010000001100111000011000;
   assign mem[90175:90144] = 32'b00000001001110101110100101110100;
   assign mem[90207:90176] = 32'b00000110001110001100001010000000;
   assign mem[90239:90208] = 32'b11111101011000100011001110101000;
   assign mem[90271:90240] = 32'b11111111011011000011010110100101;
   assign mem[90303:90272] = 32'b00000011100101110110010000001000;
   assign mem[90335:90304] = 32'b11111100110011111100100110100000;
   assign mem[90367:90336] = 32'b00000011000000001110101111011100;
   assign mem[90399:90368] = 32'b00000000110001011011000000101000;
   assign mem[90431:90400] = 32'b11111001111001101010101000001000;
   assign mem[90463:90432] = 32'b11111111010110010001011011101010;
   assign mem[90495:90464] = 32'b11111100001111001101101100001000;
   assign mem[90527:90496] = 32'b00000000000110011110110011110000;
   assign mem[90559:90528] = 32'b11110111001110010111001001000000;
   assign mem[90591:90560] = 32'b11111101111011010100010010001000;
   assign mem[90623:90592] = 32'b00000111001110001011010010110000;
   assign mem[90655:90624] = 32'b11101000010101100111000001100000;
   assign mem[90687:90656] = 32'b11100010100010010101101001000000;
   assign mem[90719:90688] = 32'b00001110101000101100111101110000;
   assign mem[90751:90720] = 32'b00001011001100101010011111110000;
   assign mem[90783:90752] = 32'b00000101100110001111000000011000;
   assign mem[90815:90784] = 32'b11111111001110000001111010110100;
   assign mem[90847:90816] = 32'b11111100011101100011000111001100;
   assign mem[90879:90848] = 32'b11110010011010001001110101100000;
   assign mem[90911:90880] = 32'b00000100011101111000100010111000;
   assign mem[90943:90912] = 32'b11111110100000110000100111001000;
   assign mem[90975:90944] = 32'b11111010010111100001100010000000;
   assign mem[91007:90976] = 32'b11111110010111101000110101001110;
   assign mem[91039:91008] = 32'b11111011010101101000010110100000;
   assign mem[91071:91040] = 32'b00000101111001101100111000010000;
   assign mem[91103:91072] = 32'b00000000011010010110010000001000;
   assign mem[91135:91104] = 32'b00000100001111101100110010011000;
   assign mem[91167:91136] = 32'b11111100011110001110010110000000;
   assign mem[91199:91168] = 32'b11111011000000010111000110100000;
   assign mem[91231:91200] = 32'b00000011101001011110001111010000;
   assign mem[91263:91232] = 32'b00000001111101110010011101111010;
   assign mem[91295:91264] = 32'b00000000100000100100100001001101;
   assign mem[91327:91296] = 32'b00000000000111011111101010011000;
   assign mem[91359:91328] = 32'b11111101000101000111110111000100;
   assign mem[91391:91360] = 32'b11111111001001000110010110000000;
   assign mem[91423:91392] = 32'b11111111000010110011001110101000;
   assign mem[91455:91424] = 32'b00000010001010111010100100100000;
   assign mem[91487:91456] = 32'b00000000010101001100101111011001;
   assign mem[91519:91488] = 32'b00000001010000000111001100110000;
   assign mem[91551:91520] = 32'b11111000001011100001010000100000;
   assign mem[91583:91552] = 32'b00000101110001101111001100100000;
   assign mem[91615:91584] = 32'b11110111110101100000111011110000;
   assign mem[91647:91616] = 32'b00000110100011001001101000011000;
   assign mem[91679:91648] = 32'b00001001100111110111111001100000;
   assign mem[91711:91680] = 32'b11111010000001100101011111101000;
   assign mem[91743:91712] = 32'b11111111111000000001111110001000;
   assign mem[91775:91744] = 32'b11111011101000101011000010110000;
   assign mem[91807:91776] = 32'b00000101110110000011011000100000;
   assign mem[91839:91808] = 32'b11111001010010010011110010101000;
   assign mem[91871:91840] = 32'b11110111101010111110110001110000;
   assign mem[91903:91872] = 32'b11110100011010100010011001110000;
   assign mem[91935:91904] = 32'b11111100001110111101010001111100;
   assign mem[91967:91936] = 32'b11110011010110010001101111010000;
   assign mem[91999:91968] = 32'b11111100001101010100001011001000;
   assign mem[92031:92000] = 32'b00001000010111100111010000110000;
   assign mem[92063:92032] = 32'b00001101100011010010011110100000;
   assign mem[92095:92064] = 32'b11110001100101101000000110100000;
   assign mem[92127:92096] = 32'b00000000100110110000011111101001;
   assign mem[92159:92128] = 32'b11111001100110001101000110001000;
   assign mem[92191:92160] = 32'b11111100011010001101100010110100;
   assign mem[92223:92192] = 32'b00001001100101111110110001010000;
   assign mem[92255:92224] = 32'b11110111001101001111110010000000;
   assign mem[92287:92256] = 32'b11111011111100100110100101101000;
   assign mem[92319:92288] = 32'b00000101111110000100000001101000;
   assign mem[92351:92320] = 32'b00000001101110000111011010011110;
   assign mem[92383:92352] = 32'b11111100000011101010100110100000;
   assign mem[92415:92384] = 32'b00000100001111111011001101001000;
   assign mem[92447:92416] = 32'b11111010110101010100010001011000;
   assign mem[92479:92448] = 32'b11111011010101101101101110010000;
   assign mem[92511:92480] = 32'b11111000101101001101001001000000;
   assign mem[92543:92512] = 32'b00001010010000101111111110110000;
   assign mem[92575:92544] = 32'b11110000010101011110000011000000;
   assign mem[92607:92576] = 32'b11110000101010000101111000100000;
   assign mem[92639:92608] = 32'b00001101000111011111110010000000;
   assign mem[92671:92640] = 32'b11111110010110110010110100001000;
   assign mem[92703:92672] = 32'b00000001001001101101101010001010;
   assign mem[92735:92704] = 32'b11110111011101000011000000110000;
   assign mem[92767:92736] = 32'b00000110000001000101001011010000;
   assign mem[92799:92768] = 32'b11110110010101000010010110000000;
   assign mem[92831:92800] = 32'b00000010110010010000010010100100;
   assign mem[92863:92832] = 32'b11111001011001110001101000011000;
   assign mem[92895:92864] = 32'b11111010100011011011001010001000;
   assign mem[92927:92896] = 32'b11111100111011110111110001111100;
   assign mem[92959:92928] = 32'b00000011010101001001000100001100;
   assign mem[92991:92960] = 32'b00001000001011111010101000010000;
   assign mem[93023:92992] = 32'b00000010001000100000000111011000;
   assign mem[93055:93024] = 32'b11110100001001111100010111010000;
   assign mem[93087:93056] = 32'b00000001000000001110000101101000;
   assign mem[93119:93088] = 32'b00000001001101100111101001101110;
   assign mem[93151:93120] = 32'b11101001110110101110011100100000;
   assign mem[93183:93152] = 32'b00000101000010101111001011010000;
   assign mem[93215:93184] = 32'b11111001001001100010000100010000;
   assign mem[93247:93216] = 32'b00001000000111101110001110100000;
   assign mem[93279:93248] = 32'b00000000000101001010111110011011;
   assign mem[93311:93280] = 32'b00001000001100001100110101100000;
   assign mem[93343:93312] = 32'b00000101101110110000100101111000;
   assign mem[93375:93344] = 32'b00000001001100101011000001111110;
   assign mem[93407:93376] = 32'b11111111110001011110010110000011;
   assign mem[93439:93408] = 32'b11110100000010001000011011110000;
   assign mem[93471:93440] = 32'b00000110110010001101001101111000;
   assign mem[93503:93472] = 32'b00000011100001101100101111001000;
   assign mem[93535:93504] = 32'b00000010011101111000001010111100;
   assign mem[93567:93536] = 32'b11111111110011010000101110111111;
   assign mem[93599:93568] = 32'b11111101000111111011111011111000;
   assign mem[93631:93600] = 32'b11111101011110011001000100000000;
   assign mem[93663:93632] = 32'b11111111110101101100111010111001;
   assign mem[93695:93664] = 32'b00000001111111000100011100110100;
   assign mem[93727:93696] = 32'b00000011011111111000010100101000;
   assign mem[93759:93728] = 32'b00000001111010111110110000111110;
   assign mem[93791:93760] = 32'b00000010011000111000101000000000;
   assign mem[93823:93792] = 32'b11111110101000010101111010001100;
   assign mem[93855:93824] = 32'b11111111001000110000101111101011;
   assign mem[93887:93856] = 32'b00000100110111010101010001001000;
   assign mem[93919:93888] = 32'b11110111000011110010001000100000;
   assign mem[93951:93920] = 32'b11111100000011001111110101101100;
   assign mem[93983:93952] = 32'b11111101001010000101111110010000;
   assign mem[94015:93984] = 32'b00000000001101111110000000111001;
   assign mem[94047:94016] = 32'b00000011000000101011010011001100;
   assign mem[94079:94048] = 32'b00000001110100111010001001100100;
   assign mem[94111:94080] = 32'b00000101001101010101010011001000;
   assign mem[94143:94112] = 32'b11111101010111001110011010001000;
   assign mem[94175:94144] = 32'b11111101001100110001110001101100;
   assign mem[94207:94176] = 32'b11111100111100100101110100011100;
   assign mem[94239:94208] = 32'b00000000110110011111010011111111;
   assign mem[94271:94240] = 32'b00000101000000010001000000100000;
   assign mem[94303:94272] = 32'b00000001010001000111110111110110;
   assign mem[94335:94304] = 32'b11111011100101110001100010001000;
   assign mem[94367:94336] = 32'b11111100011101111110110101111100;
   assign mem[94399:94368] = 32'b11111101111011000000100100101100;
   assign mem[94431:94400] = 32'b00000001000100011101111111110010;
   assign mem[94463:94432] = 32'b00000110111011001101101000010000;
   assign mem[94495:94464] = 32'b11100110110011110011101001100000;
   assign mem[94527:94496] = 32'b11101011101010101110011100100000;
   assign mem[94559:94528] = 32'b00001100100011100110001000100000;
   assign mem[94591:94560] = 32'b00010010111010000010010001000000;
   assign mem[94623:94592] = 32'b11111110100100001011110011111110;
   assign mem[94655:94624] = 32'b00000011011101010011001111100100;
   assign mem[94687:94656] = 32'b00000000001000011111011011011101;
   assign mem[94719:94688] = 32'b11101111010111010110111010100000;
   assign mem[94751:94720] = 32'b00000101011011101000101010101000;
   assign mem[94783:94752] = 32'b11111010101001111001110101101000;
   assign mem[94815:94784] = 32'b11111011010101110011110110100000;
   assign mem[94847:94816] = 32'b11111011101011011010111111110000;
   assign mem[94879:94848] = 32'b11111001011100111110110001111000;
   assign mem[94911:94880] = 32'b11111010100101110110000101011000;
   assign mem[94943:94912] = 32'b00001000000101001010110111000000;
   assign mem[94975:94944] = 32'b11111000001100010110101101111000;
   assign mem[95007:94976] = 32'b00001100100111011001001001110000;
   assign mem[95039:95008] = 32'b11111100111010010010011010111100;
   assign mem[95071:95040] = 32'b11111100011010100001101101110000;
   assign mem[95103:95072] = 32'b00000000010111001001111010000111;
   assign mem[95135:95104] = 32'b11101000011111000000001100000000;
   assign mem[95167:95136] = 32'b11101111010001000001000110100000;
   assign mem[95199:95168] = 32'b00000001100111110011010011100110;
   assign mem[95231:95200] = 32'b00001001010100011101001101000000;
   assign mem[95263:95232] = 32'b00001100001011011101010101100000;
   assign mem[95295:95264] = 32'b11111010100001110100110001110000;
   assign mem[95327:95296] = 32'b00000011001110100111110011110000;
   assign mem[95359:95328] = 32'b11110011011101000011111001010000;
   assign mem[95391:95360] = 32'b11111100011111011100111000010000;
   assign mem[95423:95392] = 32'b00001001010010101000110100110000;
   assign mem[95455:95424] = 32'b11111000110101100010100010110000;
   assign mem[95487:95456] = 32'b11111001101100101011111100101000;
   assign mem[95519:95488] = 32'b11110010110110100110001011010000;
   assign mem[95551:95520] = 32'b00000110111001001100100001011000;
   assign mem[95583:95552] = 32'b00001000011110010000011110110000;
   assign mem[95615:95584] = 32'b00000011111110001110110010001100;
   assign mem[95647:95616] = 32'b11111010110100101011110011000000;
   assign mem[95679:95648] = 32'b11111011111011101100110011111000;
   assign mem[95711:95680] = 32'b00000000010010011111100100000010;
   assign mem[95743:95712] = 32'b00000010100111011100001001110100;
   assign mem[95775:95744] = 32'b00000101110111011011001111100000;
   assign mem[95807:95776] = 32'b00000101001001100101111110000000;
   assign mem[95839:95808] = 32'b00000000011000110111011110101000;
   assign mem[95871:95840] = 32'b11111010110101010001111110011000;
   assign mem[95903:95872] = 32'b00000000010100100101111100111100;
   assign mem[95935:95904] = 32'b11111011011110101110011001110000;
   assign mem[95967:95936] = 32'b00000001001010110011110110010110;
   assign mem[95999:95968] = 32'b11111001100000111100010010111000;
   assign mem[96031:96000] = 32'b11111111100001010111010010100000;
   assign mem[96063:96032] = 32'b00000001000111010101000001010100;
   assign mem[96095:96064] = 32'b11111001101110111001000000001000;
   assign mem[96127:96096] = 32'b00000010000000110000011111100000;
   assign mem[96159:96128] = 32'b00000100011011001101010101011000;
   assign mem[96191:96160] = 32'b11111110100100001100101000011100;
   assign mem[96223:96192] = 32'b00000101001010010111100110001000;
   assign mem[96255:96224] = 32'b00000010110110111110101001001100;
   assign mem[96287:96256] = 32'b11111110000100010001111000010100;
   assign mem[96319:96288] = 32'b11111111000001111000110101101011;
   assign mem[96351:96320] = 32'b00000110100000010000111001001000;
   assign mem[96383:96352] = 32'b11111001011100101110111111000000;
   assign mem[96415:96384] = 32'b00000111101011010100111010001000;
   assign mem[96447:96416] = 32'b00000100011100110000110001011000;
   assign mem[96479:96448] = 32'b11110100000100001010010100010000;
   assign mem[96511:96480] = 32'b11110110000111110010001101100000;
   assign mem[96543:96512] = 32'b00000010011011100010101011101000;
   assign mem[96575:96544] = 32'b11111011000110011000010010101000;
   assign mem[96607:96576] = 32'b11111111010001111101111011101110;
   assign mem[96639:96608] = 32'b00000011110011100011011110000000;
   assign mem[96671:96640] = 32'b00001010110001011001001000100000;
   assign mem[96703:96672] = 32'b00000001000111100011111011000010;
   assign mem[96735:96704] = 32'b11111011000000111111011010011000;
   assign mem[96767:96736] = 32'b11110010111100110011101010100000;
   assign mem[96799:96768] = 32'b00000111001110101011101011100000;
   assign mem[96831:96800] = 32'b00000101110101010000010111010000;
   assign mem[96863:96832] = 32'b11111100001011000010000110101000;
   assign mem[96895:96864] = 32'b11111110100101000100110110001010;
   assign mem[96927:96896] = 32'b00000101101011011010110101100000;
   assign mem[96959:96928] = 32'b11101110110000100101110001000000;
   assign mem[96991:96960] = 32'b00000000011000100101111111101000;
   assign mem[97023:96992] = 32'b11111011110010100111101101110000;
   assign mem[97055:97024] = 32'b00000001011000110111001010011000;
   assign mem[97087:97056] = 32'b11111011011000100110100100111000;
   assign mem[97119:97088] = 32'b00000010010011010000011001100000;
   assign mem[97151:97120] = 32'b00000010100000010100011000011000;
   assign mem[97183:97152] = 32'b00000001010100100101101000111000;
   assign mem[97215:97184] = 32'b11111100110110011010100101001100;
   assign mem[97247:97216] = 32'b00000010110010100111011000001100;
   assign mem[97279:97248] = 32'b11111101110110101100110001010100;
   assign mem[97311:97280] = 32'b00000011010100001110010010101000;
   assign mem[97343:97312] = 32'b11111011101101001001010001011000;
   assign mem[97375:97344] = 32'b11111000111000011111100010010000;
   assign mem[97407:97376] = 32'b00000011101000111001100011001000;
   assign mem[97439:97408] = 32'b00000101101101010100111110110000;
   assign mem[97471:97440] = 32'b11111111111101100011101000010011;
   assign mem[97503:97472] = 32'b00001000010101000001000100010000;
   assign mem[97535:97504] = 32'b11111010000100101011110011001000;
   assign mem[97567:97536] = 32'b00000000101111111100001001000001;
   assign mem[97599:97568] = 32'b11111011111110010101100110011000;
   assign mem[97631:97600] = 32'b00000001010000111110100111100000;
   assign mem[97663:97632] = 32'b00001000000110000101011000010000;
   assign mem[97695:97664] = 32'b11110100010001111100011100000000;
   assign mem[97727:97696] = 32'b11110011011010001011001000000000;
   assign mem[97759:97728] = 32'b00001000100101010111011001110000;
   assign mem[97791:97760] = 32'b00001001011100100001110110110000;
   assign mem[97823:97792] = 32'b00000000100011010010101011110101;
   assign mem[97855:97824] = 32'b00000010100011010101010111100000;
   assign mem[97887:97856] = 32'b00000001110111001100001101110010;
   assign mem[97919:97888] = 32'b11111001000101000100011001110000;
   assign mem[97951:97920] = 32'b11111011101111101001011011110000;
   assign mem[97983:97952] = 32'b00000100111010110011110001111000;
   assign mem[98015:97984] = 32'b11110110011000110010101001000000;
   assign mem[98047:98016] = 32'b00000010000101000010101010011000;
   assign mem[98079:98048] = 32'b00001110101010100010011011010000;
   assign mem[98111:98080] = 32'b00000101010100100100010111001000;
   assign mem[98143:98112] = 32'b00000100011011001000000011011000;
   assign mem[98175:98144] = 32'b11111011100011111110010010000000;
   assign mem[98207:98176] = 32'b11111101001101010100111001100100;
   assign mem[98239:98208] = 32'b11111010011010101001100100011000;
   assign mem[98271:98240] = 32'b00000000100000101110110100001011;
   assign mem[98303:98272] = 32'b00001001001100100011001111010000;
   assign mem[98335:98304] = 32'b00000010011111000000011111101000;
   assign mem[98367:98336] = 32'b11111000001100100011100110000000;
   assign mem[98399:98368] = 32'b00000110111100101101111011011000;
   assign mem[98431:98400] = 32'b00000110111010000010001011100000;
   assign mem[98463:98432] = 32'b11111111100010111010001111010010;
   assign mem[98495:98464] = 32'b11111100000110111000011011010000;
   assign mem[98527:98496] = 32'b11110101001011001010000101000000;
   assign mem[98559:98528] = 32'b11110100000110110110001101110000;
   assign mem[98591:98560] = 32'b11111110111100010011101111101110;
   assign mem[98623:98592] = 32'b11110100100000001100010000000000;
   assign mem[98655:98624] = 32'b11111110100011110000010011011000;
   assign mem[98687:98656] = 32'b11111011010110110100000110100000;
   assign mem[98719:98688] = 32'b11101100011010001000110010100000;
   assign mem[98751:98720] = 32'b00001000111011101001101010100000;
   assign mem[98783:98752] = 32'b00000100001100110000000001001000;
   assign mem[98815:98784] = 32'b11110110001111001000101010110000;
   assign mem[98847:98816] = 32'b00000101110000000110110110000000;
   assign mem[98879:98848] = 32'b00000011101010101110110111010100;
   assign mem[98911:98880] = 32'b00000000111100101011100011101101;
   assign mem[98943:98912] = 32'b11110111100001000100101000110000;
   assign mem[98975:98944] = 32'b00000001111101010100001100000000;
   assign mem[99007:98976] = 32'b11111111011100100010101001010011;
   assign mem[99039:99008] = 32'b11110111001101111001001110010000;
   assign mem[99071:99040] = 32'b00000100011101011010010100100000;
   assign mem[99103:99072] = 32'b11111111010101110100011011001100;
   assign mem[99135:99104] = 32'b00000101111001001000100010010000;
   assign mem[99167:99136] = 32'b00000010010101011011001011001000;
   assign mem[99199:99168] = 32'b00000001101011111010100110100000;
   assign mem[99231:99200] = 32'b11111000010110011000110100010000;
   assign mem[99263:99232] = 32'b11111101010011101100111101000000;
   assign mem[99295:99264] = 32'b11101011100111000111011111000000;
   assign mem[99327:99296] = 32'b11111110001011011011101011100000;
   assign mem[99359:99328] = 32'b00000101111011101110000101010000;
   assign mem[99391:99360] = 32'b00000101001000001010101010111000;
   assign mem[99423:99392] = 32'b00001101100010001100111101100000;
   assign mem[99455:99424] = 32'b11110101110000101110011110000000;
   assign mem[99487:99456] = 32'b00000001010011010001010101000010;
   assign mem[99519:99488] = 32'b11111010111001011101010101111000;
   assign mem[99551:99520] = 32'b11101101111101000111010100100000;
   assign mem[99583:99552] = 32'b00000101110100010100010110010000;
   assign mem[99615:99584] = 32'b11111011101000010110110101010000;
   assign mem[99647:99616] = 32'b00000101101000010100001111110000;
   assign mem[99679:99648] = 32'b11111111100001011101100110111100;
   assign mem[99711:99680] = 32'b00000100001010011010111001110000;
   assign mem[99743:99712] = 32'b00000010000110100100111110111000;
   assign mem[99775:99744] = 32'b00000100000110101110111000001000;
   assign mem[99807:99776] = 32'b00000000001011111110111100000111;
   assign mem[99839:99808] = 32'b11110110001001100010110111100000;
   assign mem[99871:99840] = 32'b11111000011010110010111001011000;
   assign mem[99903:99872] = 32'b00000110011001010000110110000000;
   assign mem[99935:99904] = 32'b00000011011000111100010011001100;
   assign mem[99967:99936] = 32'b00001000011110110111011110010000;
   assign mem[99999:99968] = 32'b11111111101111100001110101001000;
   assign mem[100031:100000] = 32'b00000000001011111001011100000110;
   assign mem[100063:100032] = 32'b00000000111100010110010000100001;
   assign mem[100095:100064] = 32'b11110110100101110111100101110000;
   assign mem[100127:100096] = 32'b11111111101100000110010101010010;
   assign mem[100159:100128] = 32'b11111101000010010010111001010100;
   assign mem[100191:100160] = 32'b11111111001101101110000101111100;
   assign mem[100223:100192] = 32'b11110100100110011101110110000000;
   assign mem[100255:100224] = 32'b11111110010001010001100000110000;
   assign mem[100287:100256] = 32'b00000010101011111000011001101000;
   assign mem[100319:100288] = 32'b11110000000011001001100110010000;
   assign mem[100351:100320] = 32'b11110101000011000111000001010000;
   assign mem[100383:100352] = 32'b11111110111111001110111001101110;
   assign mem[100415:100384] = 32'b11110110101111010001010111100000;
   assign mem[100447:100416] = 32'b00001010001011011001101111100000;
   assign mem[100479:100448] = 32'b11110000110001010101010111010000;
   assign mem[100511:100480] = 32'b00000001000100011010011001100000;
   assign mem[100543:100512] = 32'b11111101100101011000000011011000;
   assign mem[100575:100544] = 32'b11111011111001110110001101111000;
   assign mem[100607:100576] = 32'b00000000011001100111100111011001;
   assign mem[100639:100608] = 32'b11111111011110000011000011001111;
   assign mem[100671:100640] = 32'b11111101001110001100110001001100;
   assign mem[100703:100672] = 32'b11110111101011001110111101100000;
   assign mem[100735:100704] = 32'b00000001100010010110101010001100;
   assign mem[100767:100736] = 32'b00000011010101001110101011111000;
   assign mem[100799:100768] = 32'b00000000100111000011011000011000;
   assign mem[100831:100800] = 32'b00000110000001100101111111001000;
   assign mem[100863:100832] = 32'b11111100001100001000001011110100;
   assign mem[100895:100864] = 32'b00000001111001011000001000001110;
   assign mem[100927:100896] = 32'b00000001011110111100000100001000;
   assign mem[100959:100928] = 32'b00000010000111110111010011000100;
   assign mem[100991:100960] = 32'b11111101110010011110010011101100;
   assign mem[101023:100992] = 32'b11111011001010011111111010101000;
   assign mem[101055:101024] = 32'b00000100100010001101110100011000;
   assign mem[101087:101056] = 32'b11111101101010010000110101001100;
   assign mem[101119:101088] = 32'b11111011101010000100001100011000;
   assign mem[101151:101120] = 32'b00000001110001001110110000100000;
   assign mem[101183:101152] = 32'b00000110000001101001010110110000;
   assign mem[101215:101184] = 32'b11110100010101100000010010010000;
   assign mem[101247:101216] = 32'b11110110011000001001000110000000;
   assign mem[101279:101248] = 32'b00000111101001100010100101100000;
   assign mem[101311:101280] = 32'b00001100001010000000111010010000;
   assign mem[101343:101312] = 32'b11111110111100110000101010111100;
   assign mem[101375:101344] = 32'b00000001100010011000010110110000;
   assign mem[101407:101376] = 32'b00000001110010101110001100001110;
   assign mem[101439:101408] = 32'b11111000010000110001101101011000;
   assign mem[101471:101440] = 32'b11111010001110110000111100001000;
   assign mem[101503:101472] = 32'b00000011110110110011101011111000;
   assign mem[101535:101504] = 32'b11101101110101101111110010000000;
   assign mem[101567:101536] = 32'b11110010001001001110011110000000;
   assign mem[101599:101568] = 32'b00001000111000000000001110010000;
   assign mem[101631:101600] = 32'b00000110100000100100110010111000;
   assign mem[101663:101632] = 32'b11111010001110010101001101000000;
   assign mem[101695:101664] = 32'b00000100011100001111111110101000;
   assign mem[101727:101696] = 32'b11111110011000110100101000000000;
   assign mem[101759:101728] = 32'b11111111101001010100110110110110;
   assign mem[101791:101760] = 32'b11111001110110000010010110000000;
   assign mem[101823:101792] = 32'b00001100001111011100011101000000;
   assign mem[101855:101824] = 32'b11101001001011101100010001100000;
   assign mem[101887:101856] = 32'b11101001101100001011101101100000;
   assign mem[101919:101888] = 32'b00001011010101100110100000110000;
   assign mem[101951:101920] = 32'b00000000011001000011110101001101;
   assign mem[101983:101952] = 32'b11111001001010010001100011100000;
   assign mem[102015:101984] = 32'b11111100101111100000111111111100;
   assign mem[102047:102016] = 32'b00000110010011011011011010101000;
   assign mem[102079:102048] = 32'b11101010101001111010000101100000;
   assign mem[102111:102080] = 32'b11111110111010110101000101010000;
   assign mem[102143:102112] = 32'b00000101011100110000100111001000;
   assign mem[102175:102144] = 32'b11110111101111000100001111000000;
   assign mem[102207:102176] = 32'b11110101100010001111000101000000;
   assign mem[102239:102208] = 32'b00000010100101101000101100110100;
   assign mem[102271:102240] = 32'b00001011111110110010110000100000;
   assign mem[102303:102272] = 32'b11110111111110010111111010100000;
   assign mem[102335:102304] = 32'b11111111110001110111001011100011;
   assign mem[102367:102336] = 32'b11111110001111110111011000010000;
   assign mem[102399:102368] = 32'b11111001000111100110110111101000;
   assign mem[102431:102400] = 32'b00000001010111000011011101110000;
   assign mem[102463:102432] = 32'b11111000011101111010110100010000;
   assign mem[102495:102464] = 32'b11111010000110110111000111010000;
   assign mem[102527:102496] = 32'b11111111110000110101100101100000;
   assign mem[102559:102528] = 32'b11111110011111000111011101110100;
   assign mem[102591:102560] = 32'b11111111100101110100000001001000;
   assign mem[102623:102592] = 32'b11111110010110110100111110100100;
   assign mem[102655:102624] = 32'b00000000010010111010000010100011;
   assign mem[102687:102656] = 32'b00000101000101101010100000000000;
   assign mem[102719:102688] = 32'b00000101000010000010011110111000;
   assign mem[102751:102720] = 32'b11110110101010000000110110100000;
   assign mem[102783:102752] = 32'b11111001111100111100000100110000;
   assign mem[102815:102784] = 32'b11111110101110010001101000100000;
   assign mem[102847:102816] = 32'b00000011000000001100101111010000;
   assign mem[102879:102848] = 32'b00000100011100010000010100101000;
   assign mem[102911:102880] = 32'b11111100110010101110000010000000;
   assign mem[102943:102912] = 32'b11111111110110101110111101001000;
   assign mem[102975:102944] = 32'b00001100011111011010100111010000;
   assign mem[103007:102976] = 32'b00000011011010101110011000010100;
   assign mem[103039:103008] = 32'b11111101110111000001101001100000;
   assign mem[103071:103040] = 32'b11111100011010001101000101001000;
   assign mem[103103:103072] = 32'b11111100000110010111111100111100;
   assign mem[103135:103104] = 32'b11101111101001111010111001100000;
   assign mem[103167:103136] = 32'b11110101001101110000001001010000;
   assign mem[103199:103168] = 32'b00001101111010101010111010010000;
   assign mem[103231:103200] = 32'b11111101101100100101010010100100;
   assign mem[103263:103232] = 32'b11110111110100101000011100110000;
   assign mem[103295:103264] = 32'b00001011111000011100100111010000;
   assign mem[103327:103296] = 32'b00000110101010011111001011010000;
   assign mem[103359:103328] = 32'b11110100011111000100000111000000;
   assign mem[103391:103360] = 32'b11111100011110001100011101001100;
   assign mem[103423:103392] = 32'b11111011101000011110010011000000;
   assign mem[103455:103424] = 32'b00000010000001001001110011101100;
   assign mem[103487:103456] = 32'b00000101111101001101000110011000;
   assign mem[103519:103488] = 32'b11111110101000100000011001100000;
   assign mem[103551:103520] = 32'b11111000000110110101000000000000;
   assign mem[103583:103552] = 32'b11111010010000001101011101010000;
   assign mem[103615:103584] = 32'b00000000110000111100010110111000;
   assign mem[103647:103616] = 32'b11111111001011000100110000010000;
   assign mem[103679:103648] = 32'b11110101010110001111001011010000;
   assign mem[103711:103680] = 32'b11111101101000011111010111110000;
   assign mem[103743:103712] = 32'b11111101100011111000111110101000;
   assign mem[103775:103744] = 32'b00000101100110010001101000000000;
   assign mem[103807:103776] = 32'b00001010110010110110101000110000;
   assign mem[103839:103808] = 32'b11111010100010110100001100111000;
   assign mem[103871:103840] = 32'b11110100101010100100110000110000;
   assign mem[103903:103872] = 32'b00000100001100000110110101100000;
   assign mem[103935:103904] = 32'b00000011000100110100110110001100;
   assign mem[103967:103936] = 32'b11111001110001101011011011001000;
   assign mem[103999:103968] = 32'b11110011011000101101111011110000;
   assign mem[104031:104000] = 32'b00000000101011111001010001110100;
   assign mem[104063:104032] = 32'b11111111111010010010011000100111;
   assign mem[104095:104064] = 32'b00000101010111110001110110111000;
   assign mem[104127:104096] = 32'b11110011100110001010011000000000;
   assign mem[104159:104128] = 32'b11110111000101101101010010100000;
   assign mem[104191:104160] = 32'b11111010011000011010111000110000;
   assign mem[104223:104192] = 32'b00000101000001101101011101111000;
   assign mem[104255:104224] = 32'b11111111100010010001011101111001;
   assign mem[104287:104256] = 32'b00000000110110011010000010010010;
   assign mem[104319:104288] = 32'b00001010101111100011100000100000;
   assign mem[104351:104320] = 32'b11111011001001010101001011011000;
   assign mem[104383:104352] = 32'b00000001011110100010000110100000;
   assign mem[104415:104384] = 32'b11111110101100110001110001110010;
   assign mem[104447:104416] = 32'b00000000110110010111110011100110;
   assign mem[104479:104448] = 32'b11111000100111111010111101010000;
   assign mem[104511:104480] = 32'b11111110101101111010010010111000;
   assign mem[104543:104512] = 32'b00000110000110000001110011110000;
   assign mem[104575:104544] = 32'b11111000101100100001101100011000;
   assign mem[104607:104576] = 32'b00001000010000000111000001110000;
   assign mem[104639:104608] = 32'b11111111110010111011100011000000;
   assign mem[104671:104640] = 32'b11111010101111011001111111010000;
   assign mem[104703:104672] = 32'b11101111110101010011101010100000;
   assign mem[104735:104704] = 32'b00000111010000000101110110100000;
   assign mem[104767:104736] = 32'b00000010100011101011110010110000;
   assign mem[104799:104768] = 32'b11111101010000001110100000111100;
   assign mem[104831:104800] = 32'b11101000110111011001000111100000;
   assign mem[104863:104832] = 32'b11111110111011001101111010111110;
   assign mem[104895:104864] = 32'b11111011011010100000001000011000;
   assign mem[104927:104896] = 32'b00000000000110111000100001101111;
   assign mem[104959:104928] = 32'b00000011100011010111100010011000;
   assign mem[104991:104960] = 32'b00000110000010010111100101111000;
   assign mem[105023:104992] = 32'b11111101000110001011001110000000;
   assign mem[105055:105024] = 32'b00000011011101001100001011001000;
   assign mem[105087:105056] = 32'b11111010110011100000011010011000;
   assign mem[105119:105088] = 32'b00000001100110100110001000101010;
   assign mem[105151:105120] = 32'b11101111110001101111010110000000;
   assign mem[105183:105152] = 32'b11111110010100011001000010001100;
   assign mem[105215:105184] = 32'b00001101111011001000001101110000;
   assign mem[105247:105216] = 32'b11111111011001111001000011000111;
   assign mem[105279:105248] = 32'b11111010101011110111100000110000;
   assign mem[105311:105280] = 32'b00000001101001001110100100110000;
   assign mem[105343:105312] = 32'b11111010001010000011111110001000;
   assign mem[105375:105344] = 32'b11111011011000011000001011100000;
   assign mem[105407:105376] = 32'b11111010111101100101000110110000;
   assign mem[105439:105408] = 32'b11111110110101101000001100010100;
   assign mem[105471:105440] = 32'b00000010010000000100100110000000;
   assign mem[105503:105472] = 32'b00000100010101011101001110001000;
   assign mem[105535:105504] = 32'b00000001110010111011101000010000;
   assign mem[105567:105536] = 32'b11111111000101001100000010001100;
   assign mem[105599:105568] = 32'b00000001101011000110101000111100;
   assign mem[105631:105600] = 32'b00000100011111101110000001110000;
   assign mem[105663:105632] = 32'b11111011001100000111111101010000;
   assign mem[105695:105664] = 32'b11111100110110010100011101101100;
   assign mem[105727:105696] = 32'b00000000001110000100001000111001;
   assign mem[105759:105728] = 32'b11111010011000010100110110000000;
   assign mem[105791:105760] = 32'b11111111010000101000100100101111;
   assign mem[105823:105792] = 32'b11111101000111111000101000111000;
   assign mem[105855:105824] = 32'b11111111010010110001110000001110;
   assign mem[105887:105856] = 32'b00000001000101001000000100110000;
   assign mem[105919:105888] = 32'b00000000001001001010011011100100;
   assign mem[105951:105920] = 32'b11110110110101011100101101010000;
   assign mem[105983:105952] = 32'b00000101001101110111001011010000;
   assign mem[106015:105984] = 32'b11110110111100001101101001110000;
   assign mem[106047:106016] = 32'b00000000100110010000101101100110;
   assign mem[106079:106048] = 32'b00000110011001110100000001100000;
   assign mem[106111:106080] = 32'b00000110101100011000110001110000;
   assign mem[106143:106112] = 32'b11111000101011100001100100000000;
   assign mem[106175:106144] = 32'b00000111000101110011110111000000;
   assign mem[106207:106176] = 32'b00000011001110110001101100111100;
   assign mem[106239:106208] = 32'b11110111010111011010111111110000;
   assign mem[106271:106240] = 32'b00000101111100100011111100001000;
   assign mem[106303:106272] = 32'b11111111100010010101110010101010;
   assign mem[106335:106304] = 32'b00001011010100011011011110010000;
   assign mem[106367:106336] = 32'b00000101101100111101001101001000;
   assign mem[106399:106368] = 32'b11111111111101100000010000101110;
   assign mem[106431:106400] = 32'b11101001101111010011111000100000;
   assign mem[106463:106432] = 32'b11110110110000011010100000010000;
   assign mem[106495:106464] = 32'b00001010111100011001010011000000;
   assign mem[106527:106496] = 32'b00000011111010111101110101110100;
   assign mem[106559:106528] = 32'b11111000000001010011010010001000;
   assign mem[106591:106560] = 32'b00001001001101100100011111000000;
   assign mem[106623:106592] = 32'b00000000101111100010100011101001;
   assign mem[106655:106624] = 32'b00000110101010101010101011100000;
   assign mem[106687:106656] = 32'b11111110101111101011011001000100;
   assign mem[106719:106688] = 32'b00000010000101111101010111001100;
   assign mem[106751:106720] = 32'b11110111100100100000011101010000;
   assign mem[106783:106752] = 32'b11111011111110010111110001100000;
   assign mem[106815:106784] = 32'b00001010100101101100001001010000;
   assign mem[106847:106816] = 32'b11111011111110010111010111011000;
   assign mem[106879:106848] = 32'b11110101100110111110001011000000;
   assign mem[106911:106880] = 32'b00000000010101011101111111101000;
   assign mem[106943:106912] = 32'b11111010100110111010001100100000;
   assign mem[106975:106944] = 32'b11110100010001110010100110110000;
   assign mem[107007:106976] = 32'b00000000100111101110110010000001;
   assign mem[107039:107008] = 32'b00000100000110101010100011100000;
   assign mem[107071:107040] = 32'b11111111011011110010100111001110;
   assign mem[107103:107072] = 32'b11111111000000011111111100110010;
   assign mem[107135:107104] = 32'b00000111011101010100011010001000;
   assign mem[107167:107136] = 32'b00000110111100110011010101001000;
   assign mem[107199:107168] = 32'b00000010011101111100010100101000;
   assign mem[107231:107200] = 32'b00000100000000100111001001100000;
   assign mem[107263:107232] = 32'b11111100011000011100100110111000;
   assign mem[107295:107264] = 32'b11111100011001001111111101011000;
   assign mem[107327:107296] = 32'b11111011000101010001011010010000;
   assign mem[107359:107328] = 32'b11111110010001100101110101111000;
   assign mem[107391:107360] = 32'b00000001111010000111100100101010;
   assign mem[107423:107392] = 32'b00000010101101110111010110000100;
   assign mem[107455:107424] = 32'b11111111011010101011001111000010;
   assign mem[107487:107456] = 32'b00000001100101010100101010000000;
   assign mem[107519:107488] = 32'b00000001111010110101110110100100;
   assign mem[107551:107520] = 32'b11110001100110011001111001110000;
   assign mem[107583:107552] = 32'b11111101010101010001101001111100;
   assign mem[107615:107584] = 32'b00000010110000110100110000001100;
   assign mem[107647:107616] = 32'b00000101010100000110001000110000;
   assign mem[107679:107648] = 32'b11110011101101110100010000110000;
   assign mem[107711:107680] = 32'b11101011011011001110010001100000;
   assign mem[107743:107712] = 32'b11111110001100010001101110110100;
   assign mem[107775:107744] = 32'b00000010011011111101111001010000;
   assign mem[107807:107776] = 32'b11111110011101101010100000101000;
   assign mem[107839:107808] = 32'b11111000111101101011110100111000;
   assign mem[107871:107840] = 32'b00000100110110011001000111001000;
   assign mem[107903:107872] = 32'b00000000101101101101010001011101;
   assign mem[107935:107904] = 32'b11110110111000011101110000010000;
   assign mem[107967:107936] = 32'b11111001000011110000011110010000;
   assign mem[107999:107968] = 32'b11111110110010000001101111100010;
   assign mem[108031:108000] = 32'b00000110000100000000101101111000;
   assign mem[108063:108032] = 32'b11111011010110001010011100001000;
   assign mem[108095:108064] = 32'b00000101011111111101111101011000;
   assign mem[108127:108096] = 32'b00000000100011011011111011110100;
   assign mem[108159:108128] = 32'b00000100111100111011100101001000;
   assign mem[108191:108160] = 32'b11110101110000100111100100100000;
   assign mem[108223:108192] = 32'b00000001000010110011101011001000;
   assign mem[108255:108224] = 32'b00000110110000001000100010101000;
   assign mem[108287:108256] = 32'b00000110001100010100001100111000;
   assign mem[108319:108288] = 32'b00001000110100011011000011100000;
   assign mem[108351:108320] = 32'b11110001001101000001011010010000;
   assign mem[108383:108352] = 32'b11110100111110111100010011000000;
   assign mem[108415:108384] = 32'b00000110100100011111000110010000;
   assign mem[108447:108416] = 32'b11111010110000011100100000101000;
   assign mem[108479:108448] = 32'b11110100011000100111011111000000;
   assign mem[108511:108480] = 32'b00001001000101000110001111100000;
   assign mem[108543:108512] = 32'b11111111010101111000111110000010;
   assign mem[108575:108544] = 32'b11111011111011110100101001101000;
   assign mem[108607:108576] = 32'b11111010011010110100010111110000;
   assign mem[108639:108608] = 32'b00000011111011100010010010101100;
   assign mem[108671:108640] = 32'b11110010011000000011111010010000;
   assign mem[108703:108672] = 32'b11111100100100011000110010100100;
   assign mem[108735:108704] = 32'b11111001110011100100101101110000;
   assign mem[108767:108736] = 32'b00001001101010110101001110000000;
   assign mem[108799:108768] = 32'b00000111110110010100101100010000;
   assign mem[108831:108800] = 32'b00000001110011010111011110011000;
   assign mem[108863:108832] = 32'b11111011110011001111010010010000;
   assign mem[108895:108864] = 32'b11110101101011000001000001000000;
   assign mem[108927:108896] = 32'b11110111011011100101110100010000;
   assign mem[108959:108928] = 32'b00000010100100001101101011011000;
   assign mem[108991:108960] = 32'b00000001001000001011001111011110;
   assign mem[109023:108992] = 32'b00000001110101111010010100010100;
   assign mem[109055:109024] = 32'b11111110000110111110100100111100;
   assign mem[109087:109056] = 32'b00000001010011000101001101000110;
   assign mem[109119:109088] = 32'b00000000010011111110011010001010;
   assign mem[109151:109120] = 32'b00001000000110100111011000110000;
   assign mem[109183:109152] = 32'b00000001000001000011111111101010;
   assign mem[109215:109184] = 32'b11111111100000010001001001100101;
   assign mem[109247:109216] = 32'b00001000111001000111000101000000;
   assign mem[109279:109248] = 32'b00000101001111000110100011111000;
   assign mem[109311:109280] = 32'b11101001111111100100000011100000;
   assign mem[109343:109312] = 32'b00000000101100000000010001011001;
   assign mem[109375:109344] = 32'b00000001110010110100000000000100;
   assign mem[109407:109376] = 32'b00000100100011111110100000101000;
   assign mem[109439:109408] = 32'b00000011101111010000010100001000;
   assign mem[109471:109440] = 32'b00000100011111001101111101000000;
   assign mem[109503:109472] = 32'b00000011111101110000111011001000;
   assign mem[109535:109504] = 32'b00000010100001100110100101110000;
   assign mem[109567:109536] = 32'b00000001100011011010101100011100;
   assign mem[109599:109568] = 32'b11110101111101100001000011000000;
   assign mem[109631:109600] = 32'b11111101001001101000010100100100;
   assign mem[109663:109632] = 32'b11111110011010000001001110101110;
   assign mem[109695:109664] = 32'b11111101010100110000100110100100;
   assign mem[109727:109696] = 32'b00000100110101110011101011100000;
   assign mem[109759:109728] = 32'b00001000110111100001110111100000;
   assign mem[109791:109760] = 32'b00001011010000100000111010000000;
   assign mem[109823:109792] = 32'b00000001001011101010011011010110;
   assign mem[109855:109824] = 32'b11111011101000111101000001100000;
   assign mem[109887:109856] = 32'b11110001111100001011111101010000;
   assign mem[109919:109888] = 32'b00000100011100001001111010111000;
   assign mem[109951:109920] = 32'b00000001101011111000100110111110;
   assign mem[109983:109952] = 32'b11111011010011101001101111100000;
   assign mem[110015:109984] = 32'b00000000010101110101101100111011;
   assign mem[110047:110016] = 32'b00000011011000011101111010011000;
   assign mem[110079:110048] = 32'b00000011101101010111001100100100;
   assign mem[110111:110080] = 32'b11111011011111101000111100111000;
   assign mem[110143:110112] = 32'b00000100110001111101010000111000;
   assign mem[110175:110144] = 32'b11111000000001000011010010100000;
   assign mem[110207:110176] = 32'b11110111011100000111001111100000;
   assign mem[110239:110208] = 32'b00000001000010000110111101001000;
   assign mem[110271:110240] = 32'b00000010001001011100011000110000;
   assign mem[110303:110272] = 32'b00000010100110111101000110111000;
   assign mem[110335:110304] = 32'b00000100101110111100001110100000;
   assign mem[110367:110336] = 32'b00000101011100011101100010100000;
   assign mem[110399:110368] = 32'b00000010001010001010010011101100;
   assign mem[110431:110400] = 32'b11111010010001110100111111100000;
   assign mem[110463:110432] = 32'b00001010000100000011111001110000;
   assign mem[110495:110464] = 32'b00000010100100111000010110000000;
   assign mem[110527:110496] = 32'b00000011010011000001111111011100;
   assign mem[110559:110528] = 32'b11111000100000101011001111110000;
   assign mem[110591:110560] = 32'b11111101011101010000111010010100;
   assign mem[110623:110592] = 32'b00000110110110110011110001010000;
   assign mem[110655:110624] = 32'b11101011101110011101100110000000;
   assign mem[110687:110656] = 32'b11110111101110100011101111000000;
   assign mem[110719:110688] = 32'b00000010001000101011100110000000;
   assign mem[110751:110720] = 32'b11110001001011010111110011100000;
   assign mem[110783:110752] = 32'b00000110110011001110001111101000;
   assign mem[110815:110784] = 32'b11110010001100011100111100010000;
   assign mem[110847:110816] = 32'b11111010101100000110111101001000;
   assign mem[110879:110848] = 32'b11111110010010001001110100110100;
   assign mem[110911:110880] = 32'b00001100011001011101110111100000;
   assign mem[110943:110912] = 32'b00001101110011110010110010000000;
   assign mem[110975:110944] = 32'b11111110010010111111010100001010;
   assign mem[111007:110976] = 32'b11110101100010010100110111100000;
   assign mem[111039:111008] = 32'b11110001000101011110100111010000;
   assign mem[111071:111040] = 32'b00000011010100111000010100100100;
   assign mem[111103:111072] = 32'b11111001011110010001011000011000;
   assign mem[111135:111104] = 32'b11111111101100011001011000100100;
   assign mem[111167:111136] = 32'b11111100011110001010111111110000;
   assign mem[111199:111168] = 32'b00000001001110011010000101011000;
   assign mem[111231:111200] = 32'b11111101011010110100110010010100;
   assign mem[111263:111232] = 32'b00000001110111001000100110101000;
   assign mem[111295:111264] = 32'b00000000111111101100100101101010;
   assign mem[111327:111296] = 32'b00000000010100101111010001000111;
   assign mem[111359:111328] = 32'b00000011011100000110010110111100;
   assign mem[111391:111360] = 32'b00000000010110001011100111010111;
   assign mem[111423:111392] = 32'b11111010100101110011000010011000;
   assign mem[111455:111424] = 32'b11111110111010110000111000100000;
   assign mem[111487:111456] = 32'b00000000000001001010010010100100;
   assign mem[111519:111488] = 32'b11111100010110001000111110101000;
   assign mem[111551:111520] = 32'b11111001001001001111011001101000;
   assign mem[111583:111552] = 32'b00000010101100001111111000010100;
   assign mem[111615:111584] = 32'b00000001010011101001100001111100;
   assign mem[111647:111616] = 32'b00000000000110010111100010011101;
   assign mem[111679:111648] = 32'b00000100011110111101000010100000;
   assign mem[111711:111680] = 32'b11111111101000100100001000001101;
   assign mem[111743:111712] = 32'b00000100100111011001001110100000;
   assign mem[111775:111744] = 32'b11111111100111000000011111011011;
   assign mem[111807:111776] = 32'b11111110111011110101001101010100;
   assign mem[111839:111808] = 32'b00000011111011101100011100000100;
   assign mem[111871:111840] = 32'b11110110011001000101000001000000;
   assign mem[111903:111872] = 32'b11111101011010111000110000101100;
   assign mem[111935:111904] = 32'b00000111010010101111111101000000;
   assign mem[111967:111936] = 32'b00000011011011111011000110011100;
   assign mem[111999:111968] = 32'b11111011000000100011010111011000;
   assign mem[112031:112000] = 32'b00000000010001101111011100000111;
   assign mem[112063:112032] = 32'b00000001011000110000111110100000;
   assign mem[112095:112064] = 32'b11111010100011110010111011110000;
   assign mem[112127:112096] = 32'b00000000100000011011010101111101;
   assign mem[112159:112128] = 32'b00000010011010000101000110100100;
   assign mem[112191:112160] = 32'b11110001110111001010001101010000;
   assign mem[112223:112192] = 32'b00000101111011011001000101011000;
   assign mem[112255:112224] = 32'b00000100001001000000011000000000;
   assign mem[112287:112256] = 32'b11111011110000100010010100100000;
   assign mem[112319:112288] = 32'b11111101000111110010111110001100;
   assign mem[112351:112320] = 32'b11111000110111001110011100010000;
   assign mem[112383:112352] = 32'b00000110101101000111100111100000;
   assign mem[112415:112384] = 32'b00000110001111011000100001011000;
   assign mem[112447:112416] = 32'b00000101111001001100000001101000;
   assign mem[112479:112448] = 32'b11111111101011110000001110001110;
   assign mem[112511:112480] = 32'b11110111000101101011110111100000;
   assign mem[112543:112512] = 32'b11111110001010001010010101000000;
   assign mem[112575:112544] = 32'b00000110011010111011001011001000;
   assign mem[112607:112576] = 32'b00000010100010101111010100100000;
   assign mem[112639:112608] = 32'b11110100010100011100110100110000;
   assign mem[112671:112640] = 32'b00000111001111000100001010010000;
   assign mem[112703:112672] = 32'b11111010011100011100011111111000;
   assign mem[112735:112704] = 32'b00000001001001100001100110011010;
   assign mem[112767:112736] = 32'b11111101101010111001010011000100;
   assign mem[112799:112768] = 32'b11110101111010001000110101100000;
   assign mem[112831:112800] = 32'b11111010100011000000011000010000;
   assign mem[112863:112832] = 32'b00000001101111111101000001100100;
   assign mem[112895:112864] = 32'b11111110010000101110111000000100;
   assign mem[112927:112896] = 32'b11111110101110100110111011100000;
   assign mem[112959:112928] = 32'b00001000001000100111000110110000;
   assign mem[112991:112960] = 32'b00000010111000111000100100111100;
   assign mem[113023:112992] = 32'b11110110000000100010100010000000;
   assign mem[113055:113024] = 32'b11111001010010111100010011110000;
   assign mem[113087:113056] = 32'b11111001010110000100000011101000;
   assign mem[113119:113088] = 32'b11111101101001110100000001001100;
   assign mem[113151:113120] = 32'b11111110010000011011110101100000;
   assign mem[113183:113152] = 32'b00000001010100000100111100001010;
   assign mem[113215:113184] = 32'b11111001001110100010010110010000;
   assign mem[113247:113216] = 32'b11111111011010001110010011010100;
   assign mem[113279:113248] = 32'b00001000110010001111110010110000;
   assign mem[113311:113280] = 32'b11110101101101001010000111010000;
   assign mem[113343:113312] = 32'b00000100100111011100101011110000;
   assign mem[113375:113344] = 32'b11111011001110101100011111000000;
   assign mem[113407:113376] = 32'b00000010111110011011010000110100;
   assign mem[113439:113408] = 32'b11111100110110101111010001111000;
   assign mem[113471:113440] = 32'b11110110110000101000010000110000;
   assign mem[113503:113472] = 32'b11111100000100111110010011100000;
   assign mem[113535:113504] = 32'b00000100100101001110100001100000;
   assign mem[113567:113536] = 32'b00001010001010001000000111010000;
   assign mem[113599:113568] = 32'b11110101000000110111010001100000;
   assign mem[113631:113600] = 32'b11111101000000101001001010001000;
   assign mem[113663:113632] = 32'b11111100011111000001000101110100;
   assign mem[113695:113664] = 32'b00000101000001101100001000100000;
   assign mem[113727:113696] = 32'b11111011110010001011111101100000;
   assign mem[113759:113728] = 32'b00000001001110011110110001000000;
   assign mem[113791:113760] = 32'b11111000100111011011001011010000;
   assign mem[113823:113792] = 32'b00000010100000110011110000100000;
   assign mem[113855:113824] = 32'b11111010101110010100111110110000;
   assign mem[113887:113856] = 32'b00000101101110100100001110001000;
   assign mem[113919:113888] = 32'b00000000111011000011011001100010;
   assign mem[113951:113920] = 32'b11110010101111000000110011000000;
   assign mem[113983:113952] = 32'b11111111101110000001111000110010;
   assign mem[114015:113984] = 32'b00000101111101100000111100010000;
   assign mem[114047:114016] = 32'b00000010100011010010011111111000;
   assign mem[114079:114048] = 32'b00000000101011101001110000011000;
   assign mem[114111:114080] = 32'b11101100101011001111010000000000;
   assign mem[114143:114112] = 32'b11110111100111011100000101110000;
   assign mem[114175:114144] = 32'b00010001101010111001000111000000;
   assign mem[114207:114176] = 32'b11111101111110000101010101100100;
   assign mem[114239:114208] = 32'b11110010011011101010110111100000;
   assign mem[114271:114240] = 32'b00000011101100111001011101010100;
   assign mem[114303:114272] = 32'b00000101001001101110011111110000;
   assign mem[114335:114304] = 32'b11111011001100111110011011101000;
   assign mem[114367:114336] = 32'b11110110110001110011010100010000;
   assign mem[114399:114368] = 32'b11111111010000100001001100000010;
   assign mem[114431:114400] = 32'b11111110001101000010100010101100;
   assign mem[114463:114432] = 32'b00000011011110110011100101000000;
   assign mem[114495:114464] = 32'b00001010111000111010011001110000;
   assign mem[114527:114496] = 32'b11111101101111100111100110100000;
   assign mem[114559:114528] = 32'b11111110000111101110010001101010;
   assign mem[114591:114560] = 32'b11111110000100001010011111100110;
   assign mem[114623:114592] = 32'b11110100010011111001100000010000;
   assign mem[114655:114624] = 32'b11111110101100010000001010110000;
   assign mem[114687:114656] = 32'b00000011100101000001000111001000;
   assign mem[114719:114688] = 32'b00000101010110010110010011111000;
   assign mem[114751:114720] = 32'b11111110000100110111111100010100;
   assign mem[114783:114752] = 32'b00000010100110011010110011110100;
   assign mem[114815:114784] = 32'b00001010110011111011011111000000;
   assign mem[114847:114816] = 32'b00000111100000101010000011000000;
   assign mem[114879:114848] = 32'b11110000110100010111001000100000;
   assign mem[114911:114880] = 32'b00000100110000101011001101010000;
   assign mem[114943:114912] = 32'b11110100000011111001000100000000;
   assign mem[114975:114944] = 32'b00000010111101100101110110000000;
   assign mem[115007:114976] = 32'b00000001011010100110101100111110;
   assign mem[115039:115008] = 32'b00000111010000000110110011011000;
   assign mem[115071:115040] = 32'b11110010001111101111111011100000;
   assign mem[115103:115072] = 32'b00000000110100000100110010010100;
   assign mem[115135:115104] = 32'b11111100101000010110110111101000;
   assign mem[115167:115136] = 32'b11111101010111101000001011110100;
   assign mem[115199:115168] = 32'b11111100001110100010110000000000;
   assign mem[115231:115200] = 32'b11111011011011011110111101110000;
   assign mem[115263:115232] = 32'b11111111100011101000100010010111;
   assign mem[115295:115264] = 32'b11110011101110110001101011100000;
   assign mem[115327:115296] = 32'b11111111010011111010001011011111;
   assign mem[115359:115328] = 32'b00000111000000011101101011111000;
   assign mem[115391:115360] = 32'b11111101101110111110100110110100;
   assign mem[115423:115392] = 32'b11111010111110001111011011110000;
   assign mem[115455:115424] = 32'b11111110010111000101101001101110;
   assign mem[115487:115456] = 32'b00001011000101010111010010110000;
   assign mem[115519:115488] = 32'b00000010101111100000111110001100;
   assign mem[115551:115520] = 32'b11110010111101100010111111010000;
   assign mem[115583:115552] = 32'b11110111110010001101011000010000;
   assign mem[115615:115584] = 32'b00000110110010001111100001100000;
   assign mem[115647:115616] = 32'b00000010101111100101111000100000;
   assign mem[115679:115648] = 32'b11110100010111111000001010100000;
   assign mem[115711:115680] = 32'b11110000001110000100111111110000;
   assign mem[115743:115712] = 32'b00000001111100100001000110001110;
   assign mem[115775:115744] = 32'b00000000101100010011001011110000;
   assign mem[115807:115776] = 32'b11110110101111001000011001000000;
   assign mem[115839:115808] = 32'b11110001000101100011010010100000;
   assign mem[115871:115840] = 32'b11110110001001010101110110000000;
   assign mem[115903:115872] = 32'b11111110111111110111101111000100;
   assign mem[115935:115904] = 32'b00000001011101101110001000101000;
   assign mem[115967:115936] = 32'b00000101110111010011100101011000;
   assign mem[115999:115968] = 32'b11110011110010000100110010110000;
   assign mem[116031:116000] = 32'b11110111000011101110011010010000;
   assign mem[116063:116032] = 32'b11111110001110101011001010011010;
   assign mem[116095:116064] = 32'b00000101101101100100010111100000;
   assign mem[116127:116096] = 32'b00000001000011110000110100010010;
   assign mem[116159:116128] = 32'b11111011101001011100100001111000;
   assign mem[116191:116160] = 32'b11111000100110010001100001110000;
   assign mem[116223:116192] = 32'b00000011010111010101101011010100;
   assign mem[116255:116224] = 32'b11111011001100110101000001100000;
   assign mem[116287:116256] = 32'b00000011010111000101001001001100;
   assign mem[116319:116288] = 32'b00000100101111001100001011111000;
   assign mem[116351:116320] = 32'b11111010100011100010011111100000;
   assign mem[116383:116352] = 32'b00001100111100000100101011010000;
   assign mem[116415:116384] = 32'b00000000010111010101000100110101;
   assign mem[116447:116416] = 32'b11111110100000110100011111001110;
   assign mem[116479:116448] = 32'b11111001001101000110101001111000;
   assign mem[116511:116480] = 32'b11111111111111011101001011101001;
   assign mem[116543:116512] = 32'b11111111010101011001001111100101;
   assign mem[116575:116544] = 32'b11110100011111000000111100010000;
   assign mem[116607:116576] = 32'b11111111111000110011010000000101;
   assign mem[116639:116608] = 32'b00000010110111111001111000101000;
   assign mem[116671:116640] = 32'b00000000100110111010001100011111;
   assign mem[116703:116672] = 32'b11111010110110100000111011110000;
   assign mem[116735:116704] = 32'b00000011111101010111100001001100;
   assign mem[116767:116736] = 32'b00000110010110011011001001110000;
   assign mem[116799:116768] = 32'b11111100000000110100100101000100;
   assign mem[116831:116800] = 32'b00000011010010011101011011000000;
   assign mem[116863:116832] = 32'b00000000011111100110101000110001;
   assign mem[116895:116864] = 32'b11111011010110110100110110011000;
   assign mem[116927:116896] = 32'b11111111011101011110001110011001;
   assign mem[116959:116928] = 32'b00000110111101000111000000010000;
   assign mem[116991:116960] = 32'b11111011001001001001100010110000;
   assign mem[117023:116992] = 32'b00000000101000000101001101010011;
   assign mem[117055:117024] = 32'b11111110110001111100111110110010;
   assign mem[117087:117056] = 32'b11111110000111101111000110010000;
   assign mem[117119:117088] = 32'b11111101011110101110101000100000;
   assign mem[117151:117120] = 32'b11111111111110101000011101111111;
   assign mem[117183:117152] = 32'b11111011001111000001001100111000;
   assign mem[117215:117184] = 32'b11111100010001111101100010111100;
   assign mem[117247:117216] = 32'b11111101011000010010000000011000;
   assign mem[117279:117248] = 32'b00000000101011010011011111111101;
   assign mem[117311:117280] = 32'b00000010110001111100100100100000;
   assign mem[117343:117312] = 32'b00000010100011011000100000001000;
   assign mem[117375:117344] = 32'b00000000100010101100101101010010;
   assign mem[117407:117376] = 32'b11111101011000100111101011000100;
   assign mem[117439:117408] = 32'b00000010010110001111111000011000;
   assign mem[117471:117440] = 32'b11111111100100100001000010111011;
   assign mem[117503:117472] = 32'b11111100101101100111100111100000;
   assign mem[117535:117504] = 32'b11111011101110000110111101100000;
   assign mem[117567:117536] = 32'b11111111001110101011011101011010;
   assign mem[117599:117568] = 32'b11111100010101101101000110110000;
   assign mem[117631:117600] = 32'b11111111101100011011101000001001;
   assign mem[117663:117632] = 32'b11111101111101110101100101101000;
   assign mem[117695:117664] = 32'b00000000101110111000100011101000;
   assign mem[117727:117696] = 32'b11111100110000110111001100110000;
   assign mem[117759:117728] = 32'b11111111010011101111000100010101;
   assign mem[117791:117760] = 32'b11111001100100100100011100011000;
   assign mem[117823:117792] = 32'b00000000000001110111101000101011;
   assign mem[117855:117824] = 32'b00000000010001101100101111000000;
   assign mem[117887:117856] = 32'b00000000000110110001111011100010;
   assign mem[117919:117888] = 32'b11111011110110111011101110000000;
   assign mem[117951:117920] = 32'b11111010010110001110000101100000;
   assign mem[117983:117952] = 32'b11111110101001001101110001001110;
   assign mem[118015:117984] = 32'b00000101100010001101000000000000;
   assign mem[118047:118016] = 32'b00000001001011010000010001111110;
   assign mem[118079:118048] = 32'b11110111010011110000101010000000;
   assign mem[118111:118080] = 32'b00000111110101000010100101111000;
   assign mem[118143:118112] = 32'b11111111000000000111111000001010;
   assign mem[118175:118144] = 32'b11111000111100111000111001000000;
   assign mem[118207:118176] = 32'b11111101001010000000111001001100;
   assign mem[118239:118208] = 32'b11111100100100110010111000110000;
   assign mem[118271:118240] = 32'b11111111011010010100101011110011;
   assign mem[118303:118272] = 32'b00000010111111010110110110111000;
   assign mem[118335:118304] = 32'b11111111111000010100010001100000;
   assign mem[118367:118336] = 32'b00000000101001000100010000001101;
   assign mem[118399:118368] = 32'b00000010111000001101111000101000;
   assign mem[118431:118400] = 32'b00000100101111001101110011100000;
   assign mem[118463:118432] = 32'b11111101000111100010111011111100;
   assign mem[118495:118464] = 32'b00000010011101110000110010010000;
   assign mem[118527:118496] = 32'b11111111110110011111111110010001;
   assign mem[118559:118528] = 32'b11111000000010101101001101010000;
   assign mem[118591:118560] = 32'b11111010110110110111111110101000;
   assign mem[118623:118592] = 32'b00000010101111011111110111110000;
   assign mem[118655:118624] = 32'b11111100110010111011100111110100;
   assign mem[118687:118656] = 32'b00000011000001011110011111111100;
   assign mem[118719:118688] = 32'b00001001001001010001010101100000;
   assign mem[118751:118720] = 32'b11111110010100110101101010000100;
   assign mem[118783:118752] = 32'b11111110100101110101011011000000;
   assign mem[118815:118784] = 32'b11111111100011000101001110101011;
   assign mem[118847:118816] = 32'b00000001100000001010110110001100;
   assign mem[118879:118848] = 32'b11111111010001001101101100110110;
   assign mem[118911:118880] = 32'b00000000101100011011011110101110;
   assign mem[118943:118912] = 32'b11111110111000110111001000111110;
   assign mem[118975:118944] = 32'b00000010001110100001001011111100;
   assign mem[119007:118976] = 32'b00000010100100100110001110100000;
   assign mem[119039:119008] = 32'b11111011001100101101011100011000;
   assign mem[119071:119040] = 32'b11110100010000110011010011100000;
   assign mem[119103:119072] = 32'b11111000011001001111100100001000;
   assign mem[119135:119104] = 32'b11111111010100110101110100010110;
   assign mem[119167:119136] = 32'b00000011111110010000010101011000;
   assign mem[119199:119168] = 32'b11111001101000110110111100100000;
   assign mem[119231:119200] = 32'b11111100010110100000101010010100;
   assign mem[119263:119232] = 32'b11111001111000011011000001101000;
   assign mem[119295:119264] = 32'b00000111101001101111110011100000;
   assign mem[119327:119296] = 32'b00000001010011001011001010011000;
   assign mem[119359:119328] = 32'b11111101100010101110011111101100;
   assign mem[119391:119360] = 32'b00000000100010111010001101011111;
   assign mem[119423:119392] = 32'b11111000001111000110010101110000;
   assign mem[119455:119424] = 32'b11111100000100001110001101110100;
   assign mem[119487:119456] = 32'b11111110110011100001100011000100;
   assign mem[119519:119488] = 32'b00000011101011110110101011000100;
   assign mem[119551:119520] = 32'b11110001000110011000010011010000;
   assign mem[119583:119552] = 32'b11111110000111100101100010101000;
   assign mem[119615:119584] = 32'b00000110011011010101011001011000;
   assign mem[119647:119616] = 32'b00001011110101000110011101110000;
   assign mem[119679:119648] = 32'b11111111011101101111000001111000;
   assign mem[119711:119680] = 32'b11111000110110110000111001000000;
   assign mem[119743:119712] = 32'b11111100101010101100010110010100;
   assign mem[119775:119744] = 32'b00000011011110010000011001100100;
   assign mem[119807:119776] = 32'b00000011101001000110000110001000;
   assign mem[119839:119808] = 32'b11110010101011110000110101110000;
   assign mem[119871:119840] = 32'b11111011110000000001010010011000;
   assign mem[119903:119872] = 32'b11110110010111001101011101110000;
   assign mem[119935:119904] = 32'b00000010110110111010101001001100;
   assign mem[119967:119936] = 32'b00000011000010100001100000111000;
   assign mem[119999:119968] = 32'b11111110000010011010001100110100;
   assign mem[120031:120000] = 32'b00000001100001101001111001100010;
   assign mem[120063:120032] = 32'b11111111000011100000000101110101;
   assign mem[120095:120064] = 32'b11111101011111000010000101000100;
   assign mem[120127:120096] = 32'b11111111010111001000011100001110;
   assign mem[120159:120128] = 32'b11111010100101111111011100111000;
   assign mem[120191:120160] = 32'b11111100100110010111011011011100;
   assign mem[120223:120192] = 32'b00000110110001000110110110111000;
   assign mem[120255:120224] = 32'b11111111110000100010001111010000;
   assign mem[120287:120256] = 32'b00000011111100110011100010000100;
   assign mem[120319:120288] = 32'b00000100010100000001101110101000;
   assign mem[120351:120320] = 32'b00000001101001010011001110001110;
   assign mem[120383:120352] = 32'b11111111101110010100001101010011;
   assign mem[120415:120384] = 32'b11111101011010011111001110001100;
   assign mem[120447:120416] = 32'b00000000111011001100100000001001;
   assign mem[120479:120448] = 32'b00000011000101101011010010011000;
   assign mem[120511:120480] = 32'b11111011110000100110111010101000;
   assign mem[120543:120512] = 32'b00000011110101110011010010001000;
   assign mem[120575:120544] = 32'b11111101011100101110101010000100;
   assign mem[120607:120576] = 32'b00000010011111000101000100111100;
   assign mem[120639:120608] = 32'b11111100101011111010100011101100;
   assign mem[120671:120640] = 32'b11111100101100100111010111111000;
   assign mem[120703:120672] = 32'b00000100010010110110111001111000;
   assign mem[120735:120704] = 32'b11111011100110100101111110000000;
   assign mem[120767:120736] = 32'b00000000110001010110100100101101;
   assign mem[120799:120768] = 32'b00001000010100000010111010110000;
   assign mem[120831:120800] = 32'b11111010000101111111110011010000;
   assign mem[120863:120832] = 32'b11111000000001100011101110000000;
   assign mem[120895:120864] = 32'b11111111001001110010101010000011;
   assign mem[120927:120896] = 32'b00000100100010010010110000110000;
   assign mem[120959:120928] = 32'b11111010111000010000000100101000;
   assign mem[120991:120960] = 32'b00000011110001111011101111000000;
   assign mem[121023:120992] = 32'b11111101111110010111101011010100;
   assign mem[121055:121024] = 32'b00000011111010011011100010011100;
   assign mem[121087:121056] = 32'b11111010101101101010010010000000;
   assign mem[121119:121088] = 32'b00000011110001100111110000100100;
   assign mem[121151:121120] = 32'b11110011110101101000001101000000;
   assign mem[121183:121152] = 32'b11111111011000111011111001001100;
   assign mem[121215:121184] = 32'b00000101011111100100011011111000;
   assign mem[121247:121216] = 32'b11111100001110000111001100000100;
   assign mem[121279:121248] = 32'b11111100001110001111000110111100;
   assign mem[121311:121280] = 32'b00000001011110111111011110111110;
   assign mem[121343:121312] = 32'b11111011011100110001010111000000;
   assign mem[121375:121344] = 32'b11111011100001000110101011010000;
   assign mem[121407:121376] = 32'b11111101110110011101110101100000;
   assign mem[121439:121408] = 32'b00000110000100100101000101001000;
   assign mem[121471:121440] = 32'b11111001101110010110111101010000;
   assign mem[121503:121472] = 32'b11111111101000110000100000001100;
   assign mem[121535:121504] = 32'b00000110100011110010100111010000;
   assign mem[121567:121536] = 32'b11111111111110111001010011000100;
   assign mem[121599:121568] = 32'b11111111101000100010010010001111;
   assign mem[121631:121600] = 32'b00000011101000011111000100110100;
   assign mem[121663:121632] = 32'b00000000011110011101101111000001;
   assign mem[121695:121664] = 32'b11111111000000110011010110100000;
   assign mem[121727:121696] = 32'b11111101001001101100010001010100;
   assign mem[121759:121728] = 32'b00000010010100101101111001101100;
   assign mem[121791:121760] = 32'b11110111100111010010010100100000;
   assign mem[121823:121792] = 32'b11111111100111101001010100011011;
   assign mem[121855:121824] = 32'b00000001010101011110010110110010;
   assign mem[121887:121856] = 32'b11111111011110101010110001111010;
   assign mem[121919:121888] = 32'b00000001010011110111011110011100;
   assign mem[121951:121920] = 32'b00000001101101101010111100111000;
   assign mem[121983:121952] = 32'b11111111110000111111001000011100;
   assign mem[122015:121984] = 32'b11111001010110110101101011110000;
   assign mem[122047:122016] = 32'b11111101100000110101100110010100;
   assign mem[122079:122048] = 32'b11111100001000011101010000100000;
   assign mem[122111:122080] = 32'b00000011001111011010011111101100;
   assign mem[122143:122112] = 32'b00000011001011111001110001101000;
   assign mem[122175:122144] = 32'b11111100010110101100100011111100;
   assign mem[122207:122176] = 32'b00000011100110111111000011001000;
   assign mem[122239:122208] = 32'b00000011000110100101010110101000;
   assign mem[122271:122240] = 32'b00000010011100101000011110111100;
   assign mem[122303:122272] = 32'b11111010111001110110001111110000;
   assign mem[122335:122304] = 32'b11111010101011100101100000000000;
   assign mem[122367:122336] = 32'b11111011000010111010001110000000;
   assign mem[122399:122368] = 32'b00000011101001011111111110111100;
   assign mem[122431:122400] = 32'b11111111101010011001001110001111;
   assign mem[122463:122432] = 32'b00000110101111011110011010000000;
   assign mem[122495:122464] = 32'b00000001000100110010011001111000;
   assign mem[122527:122496] = 32'b00000011001011101010110111101000;
   assign mem[122559:122528] = 32'b00000000000010111111010010110100;
   assign mem[122591:122560] = 32'b00000000100000011000000000010001;
   assign mem[122623:122592] = 32'b11110111010001010001111010000000;
   assign mem[122655:122624] = 32'b11111010110111011101000000001000;
   assign mem[122687:122656] = 32'b11111000100011111000110001011000;
   assign mem[122719:122688] = 32'b00000010111100010111111110111100;
   assign mem[122751:122720] = 32'b00000001100110010001101101101010;
   assign mem[122783:122752] = 32'b00000100011111110110100000010000;
   assign mem[122815:122784] = 32'b00000010110110001110101110001000;
   assign mem[122847:122816] = 32'b11111101001010101110101001111100;
   assign mem[122879:122848] = 32'b00000011100011000000011001111000;
   assign mem[122911:122880] = 32'b11110101001001001011111100110000;
   assign mem[122943:122912] = 32'b11111110000011110101100101000000;
   assign mem[122975:122944] = 32'b00000000111010000101101010000010;
   assign mem[123007:122976] = 32'b11111111011101110010011111010100;
   assign mem[123039:123008] = 32'b11111001110000000100011110101000;
   assign mem[123071:123040] = 32'b11111110011101000101001000001000;
   assign mem[123103:123072] = 32'b11110001011000000110101010100000;
   assign mem[123135:123104] = 32'b11111100101000101000000010110000;
   assign mem[123167:123136] = 32'b00001011101010011010010111000000;
   assign mem[123199:123168] = 32'b00001011100000101011101001000000;
   assign mem[123231:123200] = 32'b11110110001101110001110111000000;
   assign mem[123263:123232] = 32'b00000100010010110001111100110000;
   assign mem[123295:123264] = 32'b11111100101011110011001011010100;
   assign mem[123327:123296] = 32'b00000001110110100110010101000010;
   assign mem[123359:123328] = 32'b00001100011000100110100100110000;
   assign mem[123391:123360] = 32'b11111111001011100011001000100001;
   assign mem[123423:123392] = 32'b11111010110001000000110110100000;
   assign mem[123455:123424] = 32'b00001101001110111000110110100000;
   assign mem[123487:123456] = 32'b11111011101010010101010000110000;
   assign mem[123519:123488] = 32'b11100100011110100010111010100000;
   assign mem[123551:123520] = 32'b11110010010101101111011100010000;
   assign mem[123583:123552] = 32'b00000011110111000100011100000000;
   assign mem[123615:123584] = 32'b11111110001000010110011010010010;
   assign mem[123647:123616] = 32'b11110100101111110011110001010000;
   assign mem[123679:123648] = 32'b00000100010001100110110110111000;
   assign mem[123711:123680] = 32'b11111111101000010111110111010011;
   assign mem[123743:123712] = 32'b11110101010000100000010011000000;
   assign mem[123775:123744] = 32'b00000100101010111100101111110000;
   assign mem[123807:123776] = 32'b00001001101000111000000010000000;
   assign mem[123839:123808] = 32'b00001011110011011101000101010000;
   assign mem[123871:123840] = 32'b11111001111100001010011010000000;
   assign mem[123903:123872] = 32'b00000101100000001101110111100000;
   assign mem[123935:123904] = 32'b00000100000001000001011101011000;
   assign mem[123967:123936] = 32'b00000110110110110101100011011000;
   assign mem[123999:123968] = 32'b11110101000100111100110000010000;
   assign mem[124031:124000] = 32'b11111010100000110101110101111000;
   assign mem[124063:124032] = 32'b11110000011110010111001100110000;
   assign mem[124095:124064] = 32'b00000101100011100000101010000000;
   assign mem[124127:124096] = 32'b11111001000110011011000001101000;
   assign mem[124159:124128] = 32'b11110110111111010011100011000000;
   assign mem[124191:124160] = 32'b11111001000110001101001100011000;
   assign mem[124223:124192] = 32'b00000010100110001001010111110000;
   assign mem[124255:124224] = 32'b00000100100110011011100100110000;
   assign mem[124287:124256] = 32'b00001000010101001001110001100000;
   assign mem[124319:124288] = 32'b11101011101000011111100010000000;
   assign mem[124351:124320] = 32'b11110100111101011010011110100000;
   assign mem[124383:124352] = 32'b00000000010000010110010100111001;
   assign mem[124415:124384] = 32'b00000111100110101101001010000000;
   assign mem[124447:124416] = 32'b11101101000011010011010111000000;
   assign mem[124479:124448] = 32'b11111100000010011000111001000000;
   assign mem[124511:124480] = 32'b11111110010000111111010000110010;
   assign mem[124543:124512] = 32'b11110000010010100111111111100000;
   assign mem[124575:124544] = 32'b00000100000000000010011111001000;
   assign mem[124607:124576] = 32'b11110100010100100111110011000000;
   assign mem[124639:124608] = 32'b00000000001111110011000100010111;
   assign mem[124671:124640] = 32'b00000011000100100111000000100100;
   assign mem[124703:124672] = 32'b00000110001100000110010001010000;
   assign mem[124735:124704] = 32'b11111011101100001001110111011000;
   assign mem[124767:124736] = 32'b00000000101000000101110101001101;
   assign mem[124799:124768] = 32'b00000010100110110000101011011100;
   assign mem[124831:124800] = 32'b11111011001010011011111001001000;
   assign mem[124863:124832] = 32'b11111011110001001111010011101000;
   assign mem[124895:124864] = 32'b11111100000001110110100101010100;
   assign mem[124927:124896] = 32'b11101110011010000111011000100000;
   assign mem[124959:124928] = 32'b00001000101111001110101001110000;
   assign mem[124991:124960] = 32'b00000100010001101110110000000000;
   assign mem[125023:124992] = 32'b00010000100100101000001010000000;
   assign mem[125055:125024] = 32'b11101111000110010000110111100000;
   assign mem[125087:125056] = 32'b11111011111100110111101111011000;
   assign mem[125119:125088] = 32'b00000101000111010101010111110000;
   assign mem[125151:125120] = 32'b11111110000010100100010101101110;
   assign mem[125183:125152] = 32'b11111100001011101001011010101100;
   assign mem[125215:125184] = 32'b00000010110100010000010001111000;
   assign mem[125247:125216] = 32'b00001000101100110010011111110000;
   assign mem[125279:125248] = 32'b11111110010101100101011111110000;
   assign mem[125311:125280] = 32'b11111001100010100011101100001000;
   assign mem[125343:125312] = 32'b00000000010110100010001001000010;
   assign mem[125375:125344] = 32'b11111111001110000100001001001100;
   assign mem[125407:125376] = 32'b00000001000111000111000001010110;
   assign mem[125439:125408] = 32'b00000010000100010000000100001000;
   assign mem[125471:125440] = 32'b11111111011000001100010100111100;
   assign mem[125503:125472] = 32'b00000001011101100000101001111000;
   assign mem[125535:125504] = 32'b00000100001100110011000001011000;
   assign mem[125567:125536] = 32'b00000000100101011110011001101111;
   assign mem[125599:125568] = 32'b11111100101100010100011001011100;
   assign mem[125631:125600] = 32'b11111001110010010000010010001000;
   assign mem[125663:125632] = 32'b11111011111000101110011110111000;
   assign mem[125695:125664] = 32'b00001000100100100111110000110000;
   assign mem[125727:125696] = 32'b11111101011000001111000010101100;
   assign mem[125759:125728] = 32'b11110101101100100010111111010000;
   assign mem[125791:125760] = 32'b11111111011110101010001010001101;
   assign mem[125823:125792] = 32'b11111110111010000110010011010010;
   assign mem[125855:125824] = 32'b11111111001001111100101100101010;
   assign mem[125887:125856] = 32'b11110011000001001110011011100000;
   assign mem[125919:125888] = 32'b00000000000111110101111011101010;
   assign mem[125951:125920] = 32'b00000001111100101101000110111000;
   assign mem[125983:125952] = 32'b00000011101011100101000101000100;
   assign mem[126015:125984] = 32'b00000001000110011000111001000010;
   assign mem[126047:126016] = 32'b00000011000010010000001000111000;
   assign mem[126079:126048] = 32'b00000011010001101110001110110000;
   assign mem[126111:126080] = 32'b00000001101101110111001111111010;
   assign mem[126143:126112] = 32'b00000010100010111111001000100100;
   assign mem[126175:126144] = 32'b11111110100100001011111001100000;
   assign mem[126207:126176] = 32'b11111111101010101010010010110010;
   assign mem[126239:126208] = 32'b11111101100100110100000011110100;
   assign mem[126271:126240] = 32'b11111010100011010110100011101000;
   assign mem[126303:126272] = 32'b11111101110111010100111111000000;
   assign mem[126335:126304] = 32'b00000100101110001001010010100000;
   assign mem[126367:126336] = 32'b00000010110111101010000111100000;
   assign mem[126399:126368] = 32'b00000010100000110100111111100000;
   assign mem[126431:126400] = 32'b11110010010110110100010111010000;
   assign mem[126463:126432] = 32'b00000101011101010111001001100000;
   assign mem[126495:126464] = 32'b11111110000110111101111101111110;
   assign mem[126527:126496] = 32'b11111011010000100111000001110000;
   assign mem[126559:126528] = 32'b11111010101111111010010010111000;
   assign mem[126591:126560] = 32'b11111100101101100100101011111100;
   assign mem[126623:126592] = 32'b11110001111110011110111110110000;
   assign mem[126655:126624] = 32'b00000001111100011101001010100100;
   assign mem[126687:126656] = 32'b00000100100110010001101011101000;
   assign mem[126719:126688] = 32'b00000110001010011010001000001000;
   assign mem[126751:126720] = 32'b11111111101110100110010111010100;
   assign mem[126783:126752] = 32'b11111010001010101010000101001000;
   assign mem[126815:126784] = 32'b00000010101101100011001110111000;
   assign mem[126847:126816] = 32'b11110100010101100101011110000000;
   assign mem[126879:126848] = 32'b00000101101110101011110111011000;
   assign mem[126911:126880] = 32'b11111100111011101101101100100100;
   assign mem[126943:126912] = 32'b11111001010010011011001001101000;
   assign mem[126975:126944] = 32'b00000101000010000110100011011000;
   assign mem[127007:126976] = 32'b00000101101011100001001001110000;
   assign mem[127039:127008] = 32'b00000000100110101010110111001100;
   assign mem[127071:127040] = 32'b00000110000000100100001011101000;
   assign mem[127103:127072] = 32'b00000110101100010111111011110000;
   assign mem[127135:127104] = 32'b00000110111100101110000011111000;
   assign mem[127167:127136] = 32'b11110101010101101011101110100000;
   assign mem[127199:127168] = 32'b11111101000110000011101100010000;
   assign mem[127231:127200] = 32'b11111001101010011110111000111000;
   assign mem[127263:127232] = 32'b11110111001100101101110110000000;
   assign mem[127295:127264] = 32'b00001111010010010001000110100000;
   assign mem[127327:127296] = 32'b11111110101111100000101100011100;
   assign mem[127359:127328] = 32'b11110101101010010001111110100000;
   assign mem[127391:127360] = 32'b11111011110101011011100001000000;
   assign mem[127423:127392] = 32'b11111100011011100000101111011000;
   assign mem[127455:127424] = 32'b11110111110010000010011010000000;
   assign mem[127487:127456] = 32'b11110111111100101010101111110000;
   assign mem[127519:127488] = 32'b00000110101000010110101000010000;
   assign mem[127551:127520] = 32'b00000010011111100001000001010000;
   assign mem[127583:127552] = 32'b11111110011011101101011011001000;
   assign mem[127615:127584] = 32'b11111110100101110101111000101010;
   assign mem[127647:127616] = 32'b00000111100011100110100001111000;
   assign mem[127679:127648] = 32'b00001001101101101011111010110000;
   assign mem[127711:127680] = 32'b11111110001100000000000011111100;
   assign mem[127743:127712] = 32'b11111000111110110011010110111000;
   assign mem[127775:127744] = 32'b11111010011110100101100111001000;
   assign mem[127807:127776] = 32'b11111010100100100011000010111000;
   assign mem[127839:127808] = 32'b00000000011110000001011010110001;
   assign mem[127871:127840] = 32'b00000100001000110111100001111000;
   assign mem[127903:127872] = 32'b00000010100111011111101100011100;
   assign mem[127935:127904] = 32'b00000011101011111110110000001100;
   assign mem[127967:127936] = 32'b00000000100101011010000011001000;
   assign mem[127999:127968] = 32'b00000101000100101011111000101000;
   assign mem[128031:128000] = 32'b11111110110100010001010001000100;
   assign mem[128063:128032] = 32'b00000100100100110100111000100000;
   assign mem[128095:128064] = 32'b11111111010100100001110000010110;
   assign mem[128127:128096] = 32'b00000100111011111100010100100000;
   assign mem[128159:128128] = 32'b11111010110001010001100100001000;
   assign mem[128191:128160] = 32'b11111100101001001000001111010100;
   assign mem[128223:128192] = 32'b11111001110000111111100111101000;
   assign mem[128255:128224] = 32'b00000111011100110101001110000000;
   assign mem[128287:128256] = 32'b11110110010011110101011010000000;
   assign mem[128319:128288] = 32'b11111001110000001100111100000000;
   assign mem[128351:128320] = 32'b00000010111111001011011101001000;
   assign mem[128383:128352] = 32'b00000100110110011001000000110000;
   assign mem[128415:128384] = 32'b00000011101010011010001100001000;
   assign mem[128447:128416] = 32'b11110000100011110111011111100000;
   assign mem[128479:128448] = 32'b11111100010100101101111000110000;
   assign mem[128511:128480] = 32'b00000011110100101010110111110100;
   assign mem[128543:128512] = 32'b11111101100101110101011101100100;
   assign mem[128575:128544] = 32'b11111111100110000101101001011010;
   assign mem[128607:128576] = 32'b11111111101111110101110011101000;
   assign mem[128639:128608] = 32'b00000000011001111110101101101011;
   assign mem[128671:128640] = 32'b11111100110001010110100010110100;
   assign mem[128703:128672] = 32'b11110001111110001100100010010000;
   assign mem[128735:128704] = 32'b00000111001111011000101110001000;
   assign mem[128767:128736] = 32'b11110101010100001000101100000000;
   assign mem[128799:128768] = 32'b11111111010111101000101011011001;
   assign mem[128831:128800] = 32'b00000000101110001110110101101010;
   assign mem[128863:128832] = 32'b11111101100100000011001100110100;
   assign mem[128895:128864] = 32'b00000101111000101111011000001000;
   assign mem[128927:128896] = 32'b11111100010111100000101110010000;
   assign mem[128959:128928] = 32'b00001000000111010001101001000000;
   assign mem[128991:128960] = 32'b00000000001111010101101100011000;
   assign mem[129023:128992] = 32'b11111110110001100100010001010100;
   assign mem[129055:129024] = 32'b11111111001010111100111011000110;
   assign mem[129087:129056] = 32'b11111100101110100100001111001100;
   assign mem[129119:129088] = 32'b00000001000101001011100101110000;
   assign mem[129151:129120] = 32'b11110110101001001111010101000000;
   assign mem[129183:129152] = 32'b00000100011110100010001001101000;
   assign mem[129215:129184] = 32'b11111010101111000110100100001000;
   assign mem[129247:129216] = 32'b11111011110100110000100111100000;
   assign mem[129279:129248] = 32'b00000110101110100011111101011000;
   assign mem[129311:129280] = 32'b00000001000100000100101011000110;
   assign mem[129343:129312] = 32'b11111101000000101010011000001000;
   assign mem[129375:129344] = 32'b11111111100000001011111010101100;
   assign mem[129407:129376] = 32'b11110011000111101111110011100000;
   assign mem[129439:129408] = 32'b00000001111000111001110010000100;
   assign mem[129471:129440] = 32'b00000001110111101010001010101010;
   assign mem[129503:129472] = 32'b00000100100110010110100110111000;
   assign mem[129535:129504] = 32'b00000011001100010000011111101100;
   assign mem[129567:129536] = 32'b00000000111001001101111101100011;
   assign mem[129599:129568] = 32'b00000001101110111110010111001000;
   assign mem[129631:129600] = 32'b11111111100011001110101011000010;
   assign mem[129663:129632] = 32'b11111111111110110010100101111101;
   assign mem[129695:129664] = 32'b11111010010001000010111101001000;
   assign mem[129727:129696] = 32'b00000011100011110011011111101000;
   assign mem[129759:129728] = 32'b11111110101001001101011011011100;
   assign mem[129791:129760] = 32'b11111110110001011000001011001100;
   assign mem[129823:129792] = 32'b11111101110011100000101101011000;
   assign mem[129855:129824] = 32'b00000011101001011010010011100100;
   assign mem[129887:129856] = 32'b11111101011111101010110111010100;
   assign mem[129919:129888] = 32'b00000010110010010111010111010000;
   assign mem[129951:129920] = 32'b11111110001001001010100100101100;
   assign mem[129983:129952] = 32'b11111000111101001010110000100000;
   assign mem[130015:129984] = 32'b11111111011100011101110100111100;
   assign mem[130047:130016] = 32'b00000011111000101110001010001000;
   assign mem[130079:130048] = 32'b00000010101100011101001100001000;
   assign mem[130111:130080] = 32'b11111100011100011111011010101100;
   assign mem[130143:130112] = 32'b00000101000011011110001000110000;
   assign mem[130175:130144] = 32'b11111101101000100101001101110100;
   assign mem[130207:130176] = 32'b00000100110110100101110000001000;
   assign mem[130239:130208] = 32'b00000001010101100010100100001000;
   assign mem[130271:130240] = 32'b00000001011111111011111110110010;
   assign mem[130303:130272] = 32'b00000001000011100110111101001000;
   assign mem[130335:130304] = 32'b11111101111110111100001110100000;
   assign mem[130367:130336] = 32'b11101111011010101001011111000000;
   assign mem[130399:130368] = 32'b00000110110111000101001100111000;
   assign mem[130431:130400] = 32'b00000000010000000100101010010100;
   assign mem[130463:130432] = 32'b11111110000010010001011110011000;
   assign mem[130495:130464] = 32'b00000001110001001000011110101000;
   assign mem[130527:130496] = 32'b00000011100101000110100000001000;
   assign mem[130559:130528] = 32'b00000101101011101000111101101000;
   assign mem[130591:130560] = 32'b11111001111000011010111100110000;
   assign mem[130623:130592] = 32'b00000010010100100100100001000100;
   assign mem[130655:130624] = 32'b11110101001101001001000001100000;
   assign mem[130687:130656] = 32'b11110000011101111011001101010000;
   assign mem[130719:130688] = 32'b00000111110100010011000110011000;
   assign mem[130751:130720] = 32'b00000010000100110111010110110000;
   assign mem[130783:130752] = 32'b11111110011000111110110001101110;
   assign mem[130815:130784] = 32'b00000100111010001101100000100000;
   assign mem[130847:130816] = 32'b00000001010100011110010011001010;
   assign mem[130879:130848] = 32'b00000100010000001011100101111000;
   assign mem[130911:130880] = 32'b11111101101001001110010011111100;
   assign mem[130943:130912] = 32'b11111110011110101011111100001010;
   assign mem[130975:130944] = 32'b11111111010010001101100110111000;
   assign mem[131007:130976] = 32'b11111000011100010110110111111000;
   assign mem[131039:131008] = 32'b00000110010010100111001110100000;
   assign mem[131071:131040] = 32'b11111010000011111000010001110000;
   assign mem[131103:131072] = 32'b00001111010010010111101011100000;
   assign mem[131135:131104] = 32'b11110100100101101010001001100000;
   assign mem[131167:131136] = 32'b11111101010011101110001111010000;
   assign mem[131199:131168] = 32'b11111111000100011010001111101110;
   assign mem[131231:131200] = 32'b11111110101100100110100000111010;
   assign mem[131263:131232] = 32'b11111000101000100110100100010000;
   assign mem[131295:131264] = 32'b11110100110101100011101010000000;
   assign mem[131327:131296] = 32'b11100110110110011101101101100000;
   assign mem[131359:131328] = 32'b00001011100000010010111110110000;
   assign mem[131391:131360] = 32'b00000000111000000100010111010110;
   assign mem[131423:131392] = 32'b00001100010100101100011111010000;
   assign mem[131455:131424] = 32'b11111001100100011101110110110000;
   assign mem[131487:131456] = 32'b11111111000101011011110100001001;
   assign mem[131519:131488] = 32'b00000010011110011100001110000100;
   assign mem[131551:131520] = 32'b00000010100111110001110100101100;
   assign mem[131583:131552] = 32'b11111011000011000011111010010000;
   assign mem[131615:131584] = 32'b11111110001001101110101110110000;
   assign mem[131647:131616] = 32'b11111110100000000010111010000010;
   assign mem[131679:131648] = 32'b00000001101001101001000001100110;
   assign mem[131711:131680] = 32'b00000001001101100110110000010110;
   assign mem[131743:131712] = 32'b00000011110010100110100110000100;
   assign mem[131775:131744] = 32'b11111100110000101100111110111100;
   assign mem[131807:131776] = 32'b00000010011011111100010100111000;
   assign mem[131839:131808] = 32'b00000010001000111000011011010100;
   assign mem[131871:131840] = 32'b11111101100010100101011011101100;
   assign mem[131903:131872] = 32'b00000000011011101001110101011100;
   assign mem[131935:131904] = 32'b11110111010100111110011000010000;
   assign mem[131967:131936] = 32'b11111100110101010101100011001000;
   assign mem[131999:131968] = 32'b00000010111011100011011110101100;
   assign mem[132031:132000] = 32'b11111101011001111100100101101000;
   assign mem[132063:132032] = 32'b00001001011000010111101010100000;
   assign mem[132095:132064] = 32'b00000010110000110000100011000100;
   assign mem[132127:132096] = 32'b00000101011110101101100100000000;
   assign mem[132159:132128] = 32'b00000111100010001111101110001000;
   assign mem[132191:132160] = 32'b00000101000111000000110011101000;
   assign mem[132223:132192] = 32'b11111111111101011100010111010101;
   assign mem[132255:132224] = 32'b00000011010010000101001110111100;
   assign mem[132287:132256] = 32'b00000000001110011011001100101001;
   assign mem[132319:132288] = 32'b11110101100101000111011111010000;
   assign mem[132351:132320] = 32'b11111100010111110101110001101000;
   assign mem[132383:132352] = 32'b11110110000101101010111100000000;
   assign mem[132415:132384] = 32'b00000111110010101001010010000000;
   assign mem[132447:132416] = 32'b11111100001111101001001111000000;
   assign mem[132479:132448] = 32'b11111110001100101110100110110110;
   assign mem[132511:132480] = 32'b00000100111010111110010001000000;
   assign mem[132543:132512] = 32'b11101000100110111000010000100000;
   assign mem[132575:132544] = 32'b00000000100010110000101011001100;
   assign mem[132607:132576] = 32'b11111000100001101011100111101000;
   assign mem[132639:132608] = 32'b00000110111001111110101011111000;
   assign mem[132671:132640] = 32'b00000010011010101011111010001100;
   assign mem[132703:132672] = 32'b00000011111100111001001111001100;
   assign mem[132735:132704] = 32'b00000101110101111110100011010000;
   assign mem[132767:132736] = 32'b11111100100000110010101000011100;
   assign mem[132799:132768] = 32'b11111110010000000010000111001010;
   assign mem[132831:132800] = 32'b11111111111000000100000011101111;
   assign mem[132863:132832] = 32'b00000011011101100010011001111000;
   assign mem[132895:132864] = 32'b00000011111001010110010010010100;
   assign mem[132927:132896] = 32'b00000101001001001000001101111000;
   assign mem[132959:132928] = 32'b11110011001011010101111111110000;
   assign mem[132991:132960] = 32'b00000001001001011101001100101110;
   assign mem[133023:132992] = 32'b11110101101010001100110101100000;
   assign mem[133055:133024] = 32'b00000101011010101111010111000000;
   assign mem[133087:133056] = 32'b11111011011000101010100000000000;
   assign mem[133119:133088] = 32'b00000100001110001010000101000000;
   assign mem[133151:133120] = 32'b00000000001010111000011011001111;
   assign mem[133183:133152] = 32'b11110011100001010011101100110000;
   assign mem[133215:133184] = 32'b00000010110011101100111101000100;
   assign mem[133247:133216] = 32'b11111100101100010110101010010100;
   assign mem[133279:133248] = 32'b11111110011000011001001000110110;
   assign mem[133311:133280] = 32'b11111100011000100111011011011000;
   assign mem[133343:133312] = 32'b11111101011001101100100011100000;
   assign mem[133375:133344] = 32'b11111100101101001010001000101100;
   assign mem[133407:133376] = 32'b00000001000110110010001100011100;
   assign mem[133439:133408] = 32'b00000100101110100011111100101000;
   assign mem[133471:133440] = 32'b00000010000010101001000101000000;
   assign mem[133503:133472] = 32'b11111000100100001001010111000000;
   assign mem[133535:133504] = 32'b00000000010111100100100101100111;
   assign mem[133567:133536] = 32'b11111011011010010010100011111000;
   assign mem[133599:133568] = 32'b00000001000110111010101100110110;
   assign mem[133631:133600] = 32'b11111100101001100010011010011100;
   assign mem[133663:133632] = 32'b00000101001010100011000001101000;
   assign mem[133695:133664] = 32'b00000000111000011111110100101111;
   assign mem[133727:133696] = 32'b00000011001100110000101101001000;
   assign mem[133759:133728] = 32'b00000011001110011110000011101000;
   assign mem[133791:133760] = 32'b00000011100000010111100001100100;
   assign mem[133823:133792] = 32'b00000000011001101100110010000010;
   assign mem[133855:133824] = 32'b11111111000100101001010100000010;
   assign mem[133887:133856] = 32'b11111101101110010111101110110100;
   assign mem[133919:133888] = 32'b11110110001010011111001010010000;
   assign mem[133951:133920] = 32'b11111100000011000000100100010100;
   assign mem[133983:133952] = 32'b11111011110011110011001100011000;
   assign mem[134015:133984] = 32'b00000111101001101010111110001000;
   assign mem[134047:134016] = 32'b00000000010110111111111111011001;
   assign mem[134079:134048] = 32'b00001001111110100011101001000000;
   assign mem[134111:134080] = 32'b00000000111111000101011110110100;
   assign mem[134143:134112] = 32'b11111010001011100100010110101000;
   assign mem[134175:134144] = 32'b11111111110110011100100111101111;
   assign mem[134207:134176] = 32'b11111111001010011001011000111011;
   assign mem[134239:134208] = 32'b00000011000010011001000011110100;
   assign mem[134271:134240] = 32'b00000001000010001101010111100100;
   assign mem[134303:134272] = 32'b00000101111000111100110101110000;
   assign mem[134335:134304] = 32'b11111000000110000101010111000000;
   assign mem[134367:134336] = 32'b11111100110101010001101101011100;
   assign mem[134399:134368] = 32'b00000100111000100011111000011000;
   assign mem[134431:134400] = 32'b11110011111101100010100000100000;
   assign mem[134463:134432] = 32'b11111000001110100011100111110000;
   assign mem[134495:134464] = 32'b00000111000111000110111001011000;
   assign mem[134527:134496] = 32'b11111100101100101100000000110100;
   assign mem[134559:134528] = 32'b00000000101010101011000110101101;
   assign mem[134591:134560] = 32'b11111011101001000111101111010000;
   assign mem[134623:134592] = 32'b11110101011010011001010111000000;
   assign mem[134655:134624] = 32'b00001101000010110011001100010000;
   assign mem[134687:134656] = 32'b00000110010001000110110101001000;
   assign mem[134719:134688] = 32'b11111001011100101010110010011000;
   assign mem[134751:134720] = 32'b00000101011111001010011101001000;
   assign mem[134783:134752] = 32'b11111100111010010000010011111000;
   assign mem[134815:134784] = 32'b11111000011011000101011001100000;
   assign mem[134847:134816] = 32'b00000000001100100001001001010010;
   assign mem[134879:134848] = 32'b00000010110111000001011010000000;
   assign mem[134911:134880] = 32'b00000000101101110100111010001110;
   assign mem[134943:134912] = 32'b11111011111101110111001100011000;
   assign mem[134975:134944] = 32'b00001001000010010110000101100000;
   assign mem[135007:134976] = 32'b00000110001000010000001001011000;
   assign mem[135039:135008] = 32'b11110011110110001110100100110000;
   assign mem[135071:135040] = 32'b00000001010011101101110001100100;
   assign mem[135103:135072] = 32'b11111101011101010010111100111000;
   assign mem[135135:135104] = 32'b11110111011000100111100101000000;
   assign mem[135167:135136] = 32'b11111101010111001110100101001000;
   assign mem[135199:135168] = 32'b00000011100010010011100110111100;
   assign mem[135231:135200] = 32'b00000010111001100100010001110100;
   assign mem[135263:135232] = 32'b11111011111010100100100110101000;
   assign mem[135295:135264] = 32'b00000101011000011110001011000000;
   assign mem[135327:135296] = 32'b00000001111111000000000001000010;
   assign mem[135359:135328] = 32'b11111010011010111010011000001000;
   assign mem[135391:135360] = 32'b11111111011110110001001000000110;
   assign mem[135423:135392] = 32'b11111100100011100101110011101100;
   assign mem[135455:135424] = 32'b00000011111101111110110101010100;
   assign mem[135487:135456] = 32'b00001000000001101111001100110000;
   assign mem[135519:135488] = 32'b11111011111011100011101001101000;
   assign mem[135551:135520] = 32'b11111100111100100100000110011000;
   assign mem[135583:135552] = 32'b00000000000101011010110110000010;
   assign mem[135615:135584] = 32'b00000011001110110111000100111000;
   assign mem[135647:135616] = 32'b11111010011000101010101110111000;
   assign mem[135679:135648] = 32'b11111001001001100111000000010000;
   assign mem[135711:135680] = 32'b11111001100011011100111111000000;
   assign mem[135743:135712] = 32'b00000100001111001100111010100000;
   assign mem[135775:135744] = 32'b00000010100111000001111111001100;
   assign mem[135807:135776] = 32'b11110111100110000100111001110000;
   assign mem[135839:135808] = 32'b11111001110001101110100001100000;
   assign mem[135871:135840] = 32'b00000010100101110011110100111100;
   assign mem[135903:135872] = 32'b11110111000110000010001100010000;
   assign mem[135935:135904] = 32'b11111101001101000111110101000000;
   assign mem[135967:135936] = 32'b00000000110000010100101101101100;
   assign mem[135999:135968] = 32'b00001110100111110000110100100000;
   assign mem[136031:136000] = 32'b00000110011110011001100101010000;
   assign mem[136063:136032] = 32'b11111011000101100000100111110000;
   assign mem[136095:136064] = 32'b00000110001001011111110000111000;
   assign mem[136127:136096] = 32'b00000010011111111001111101011000;
   assign mem[136159:136128] = 32'b11110011100100001010010111000000;
   assign mem[136191:136160] = 32'b11111011100110000111000110111000;
   assign mem[136223:136192] = 32'b11111111010010010011100010001111;
   assign mem[136255:136224] = 32'b00000101111110101000101000010000;
   assign mem[136287:136256] = 32'b11110110110110101110101010000000;
   assign mem[136319:136288] = 32'b11111011111011010101011011010000;
   assign mem[136351:136320] = 32'b11111010001011010110111100010000;
   assign mem[136383:136352] = 32'b00000100101010010111011110100000;
   assign mem[136415:136384] = 32'b00000011110011110100101110011100;
   assign mem[136447:136416] = 32'b00001000100101100101001111010000;
   assign mem[136479:136448] = 32'b11101001110010001111011001000000;
   assign mem[136511:136480] = 32'b11111011000010100110000100110000;
   assign mem[136543:136512] = 32'b11110110100101111010001110100000;
   assign mem[136575:136544] = 32'b00000101111100111010011101100000;
   assign mem[136607:136576] = 32'b00000000001101001110011110111101;
   assign mem[136639:136608] = 32'b00000000010010000101001010001111;
   assign mem[136671:136640] = 32'b11111110011011100000010000011000;
   assign mem[136703:136672] = 32'b11111011111100010101000010111000;
   assign mem[136735:136704] = 32'b11101010100011110010011001000000;
   assign mem[136767:136736] = 32'b11110100101110110101111001000000;
   assign mem[136799:136768] = 32'b00010001011001010011001110000000;
   assign mem[136831:136800] = 32'b11111110011111110100100100100100;
   assign mem[136863:136832] = 32'b00000010001111101101110011101100;
   assign mem[136895:136864] = 32'b00001011111110100011100100100000;
   assign mem[136927:136896] = 32'b11110111011000010100100011110000;
   assign mem[136959:136928] = 32'b11110110111101100101101111010000;
   assign mem[136991:136960] = 32'b11111111101011011001101101111000;
   assign mem[137023:136992] = 32'b11111100000000100100110001100100;
   assign mem[137055:137024] = 32'b11111101000100100100110011101000;
   assign mem[137087:137056] = 32'b11110011000011000101100011010000;
   assign mem[137119:137088] = 32'b00000011100001011011011001111100;
   assign mem[137151:137120] = 32'b00000001110101110000100110011110;
   assign mem[137183:137152] = 32'b00000000011000011001011010010111;
   assign mem[137215:137184] = 32'b11111100011000110010000100100000;
   assign mem[137247:137216] = 32'b00000011110000000001100011100100;
   assign mem[137279:137248] = 32'b00001010000000010101000101100000;
   assign mem[137311:137280] = 32'b00000010011001010101010000100100;
   assign mem[137343:137312] = 32'b11111011111001011011010001000000;
   assign mem[137375:137344] = 32'b11111101001101111001000000011000;
   assign mem[137407:137376] = 32'b11111100010010011000111001011100;
   assign mem[137439:137408] = 32'b00001000100110001000001101100000;
   assign mem[137471:137440] = 32'b11110110110111100101010110110000;
   assign mem[137503:137472] = 32'b11111100011101101100111000100000;
   assign mem[137535:137504] = 32'b00001110011011100111100011010000;
   assign mem[137567:137536] = 32'b00000100101000110011011000100000;
   assign mem[137599:137568] = 32'b11111000000100011011100100111000;
   assign mem[137631:137600] = 32'b11111100001100001001011100000100;
   assign mem[137663:137632] = 32'b11111100010010101010011101000000;
   assign mem[137695:137664] = 32'b00000000011101000110110111101001;
   assign mem[137727:137696] = 32'b11111100111101100001100110000000;
   assign mem[137759:137728] = 32'b11111110010010011010000011101010;
   assign mem[137791:137760] = 32'b00000011001011110110001000101000;
   assign mem[137823:137792] = 32'b00000001110011010010111001110110;
   assign mem[137855:137824] = 32'b11111111111000100001111101001101;
   assign mem[137887:137856] = 32'b00000001010100111011001000101110;
   assign mem[137919:137888] = 32'b00000000010011001001010010001010;
   assign mem[137951:137920] = 32'b11111111010111100110010101000111;
   assign mem[137983:137952] = 32'b00000011011010100110101100000000;
   assign mem[138015:137984] = 32'b11111110011011000111010000000110;
   assign mem[138047:138016] = 32'b00000011010001100001111101101000;
   assign mem[138079:138048] = 32'b11111101010001011000101111011100;
   assign mem[138111:138080] = 32'b11111100001111011101110010101100;
   assign mem[138143:138112] = 32'b11111100111001110101000000110100;
   assign mem[138175:138144] = 32'b00000000100101111010101110010101;
   assign mem[138207:138176] = 32'b11111110111010110010110001000000;
   assign mem[138239:138208] = 32'b11111100110010101011101011100000;
   assign mem[138271:138240] = 32'b00001100011111111100100010100000;
   assign mem[138303:138272] = 32'b11110111010011000110001001100000;
   assign mem[138335:138304] = 32'b00000001100110110111010111100100;
   assign mem[138367:138336] = 32'b00000000000100111101010111001001;
   assign mem[138399:138368] = 32'b11110111001100100110110111010000;
   assign mem[138431:138400] = 32'b00000010110110011010101000000100;
   assign mem[138463:138432] = 32'b00000010011110010001000000010100;
   assign mem[138495:138464] = 32'b00000010111011011111000101000100;
   assign mem[138527:138496] = 32'b00000011011110111100100000111000;
   assign mem[138559:138528] = 32'b11111110000000110001011010100100;
   assign mem[138591:138560] = 32'b00000001111101000000010100001100;
   assign mem[138623:138592] = 32'b11111100000001001001011000000100;
   assign mem[138655:138624] = 32'b11111100011011101100100110110000;
   assign mem[138687:138656] = 32'b11111011001110101001011100001000;
   assign mem[138719:138688] = 32'b00000100001000111100100110011000;
   assign mem[138751:138720] = 32'b11111111100100010110100100100100;
   assign mem[138783:138752] = 32'b00000010111011011100111110110000;
   assign mem[138815:138784] = 32'b00000001100010010011100101000010;
   assign mem[138847:138816] = 32'b00000001000001001111000111100000;
   assign mem[138879:138848] = 32'b00000010101100001100111011000100;
   assign mem[138911:138880] = 32'b00000000110100000010110001011111;
   assign mem[138943:138912] = 32'b11111111110010000110100111001010;
   assign mem[138975:138944] = 32'b11111001111100011010110100101000;
   assign mem[139007:138976] = 32'b00000001000111010100100110011000;
   assign mem[139039:139008] = 32'b00000011011100111010010101000000;
   assign mem[139071:139040] = 32'b11111010001100010111010111010000;
   assign mem[139103:139072] = 32'b00000001101101110001110010111100;
   assign mem[139135:139104] = 32'b11111110000010100100000111001010;
   assign mem[139167:139136] = 32'b00000010000011010111010100101100;
   assign mem[139199:139168] = 32'b00000101010000100010100101000000;
   assign mem[139231:139200] = 32'b11111010000011001001011000010000;
   assign mem[139263:139232] = 32'b00000000101101010100000000010011;
   assign mem[139295:139264] = 32'b00000010001010100011111111001100;
   assign mem[139327:139296] = 32'b11111111110010011001011100110101;
   assign mem[139359:139328] = 32'b11111111101100010100110110011100;
   assign mem[139391:139360] = 32'b00000000110100110001101011011111;
   assign mem[139423:139392] = 32'b11110100111011000001111001110000;
   assign mem[139455:139424] = 32'b00000001110000000100111100111100;
   assign mem[139487:139456] = 32'b00000010000111110000110001011100;
   assign mem[139519:139488] = 32'b11111111001000111111001111111010;
   assign mem[139551:139520] = 32'b00000010111101011001101101010000;
   assign mem[139583:139552] = 32'b00000001000000111100001110000110;
   assign mem[139615:139584] = 32'b00000011001001010001000110011000;
   assign mem[139647:139616] = 32'b00000100100000010001110001110000;
   assign mem[139679:139648] = 32'b11110111111011001110101100100000;
   assign mem[139711:139680] = 32'b11111101000010010010011001111000;
   assign mem[139743:139712] = 32'b11110100111010111100011101110000;
   assign mem[139775:139744] = 32'b00000010000000101011111100000000;
   assign mem[139807:139776] = 32'b11111100001010101111001101111100;
   assign mem[139839:139808] = 32'b00000001110000001111101010010000;
   assign mem[139871:139840] = 32'b00000000010011010111010010100100;
   assign mem[139903:139872] = 32'b11110110101100110111111010010000;
   assign mem[139935:139904] = 32'b00000011001110000001000011111100;
   assign mem[139967:139936] = 32'b11111101111010100001000001011100;
   assign mem[139999:139968] = 32'b11110111001011010100001111110000;
   assign mem[140031:140000] = 32'b00000000110101010101110100010010;
   assign mem[140063:140032] = 32'b11111000100000001001110100011000;
   assign mem[140095:140064] = 32'b00000101001001110100000011111000;
   assign mem[140127:140096] = 32'b00000010001110001000100011001000;
   assign mem[140159:140128] = 32'b00001000100010101011110000000000;
   assign mem[140191:140160] = 32'b11111110011110001000010001111110;
   assign mem[140223:140192] = 32'b11111011110010111001000110000000;
   assign mem[140255:140224] = 32'b00000010010001101101110010000100;
   assign mem[140287:140256] = 32'b00000010101111100000000011010100;
   assign mem[140319:140288] = 32'b11111010101100011101101111100000;
   assign mem[140351:140320] = 32'b11111100001011110100100001101100;
   assign mem[140383:140352] = 32'b11110110111100111011010011000000;
   assign mem[140415:140384] = 32'b00000010100100010000011101000000;
   assign mem[140447:140416] = 32'b11111010101011100101011011110000;
   assign mem[140479:140448] = 32'b00000010000011111100111110011100;
   assign mem[140511:140480] = 32'b00000001011011001011110100101010;
   assign mem[140543:140512] = 32'b11110011010011110011001011110000;
   assign mem[140575:140544] = 32'b11111101111100101111100011001000;
   assign mem[140607:140576] = 32'b11111101001001001100111100101000;
   assign mem[140639:140608] = 32'b00000011100110110001010101001000;
   assign mem[140671:140640] = 32'b00000000110001000111010000011100;
   assign mem[140703:140672] = 32'b00001000101011100100010000100000;
   assign mem[140735:140704] = 32'b11110111111000101011111110110000;
   assign mem[140767:140736] = 32'b11111011000001001101000001100000;
   assign mem[140799:140768] = 32'b00000111101000110011111000101000;
   assign mem[140831:140800] = 32'b00000000110111010101001001011000;
   assign mem[140863:140832] = 32'b11111110100000111100011100111100;
   assign mem[140895:140864] = 32'b11111101111000010001110101010100;
   assign mem[140927:140896] = 32'b00000101011010011001110000011000;
   assign mem[140959:140928] = 32'b00001010010111010000000101100000;
   assign mem[140991:140960] = 32'b11111110011100110000100111110110;
   assign mem[141023:140992] = 32'b00000000011010100001010110000010;
   assign mem[141055:141024] = 32'b00000100101101001111100101001000;
   assign mem[141087:141056] = 32'b11111110100100101001111001111000;
   assign mem[141119:141088] = 32'b11101111110101011100110110000000;
   assign mem[141151:141120] = 32'b11110110110001001101110111010000;
   assign mem[141183:141152] = 32'b00000010110010010111111000111000;
   assign mem[141215:141184] = 32'b11111111001100100010011110011100;
   assign mem[141247:141216] = 32'b00000011100110110101111101011000;
   assign mem[141279:141248] = 32'b11111101111110010001000110101100;
   assign mem[141311:141280] = 32'b00000110011101010000100100100000;
   assign mem[141343:141312] = 32'b11101111110011110010010001000000;
   assign mem[141375:141344] = 32'b00000100000000001001010001101000;
   assign mem[141407:141376] = 32'b00000010100111000111000110110000;
   assign mem[141439:141408] = 32'b11111000001011100111110011110000;
   assign mem[141471:141440] = 32'b00000011100000000110010101011100;
   assign mem[141503:141472] = 32'b00000010010101010100010101001000;
   assign mem[141535:141504] = 32'b11111101010000000110011000111000;
   assign mem[141567:141536] = 32'b11111101100111011110010010000000;
   assign mem[141599:141568] = 32'b00000010111001001111110011101000;
   assign mem[141631:141600] = 32'b11111110010100010001010011111010;
   assign mem[141663:141632] = 32'b11111110110011011001001100010110;
   assign mem[141695:141664] = 32'b00001111001010100110101000010000;
   assign mem[141727:141696] = 32'b11111011000110011101001000011000;
   assign mem[141759:141728] = 32'b11110010111011010110110011000000;
   assign mem[141791:141760] = 32'b00000001111100100111100000000110;
   assign mem[141823:141792] = 32'b11111011111001001001110101100000;
   assign mem[141855:141824] = 32'b11111101000110000011001011101000;
   assign mem[141887:141856] = 32'b11111000001101001100111000100000;
   assign mem[141919:141888] = 32'b00001001000100001111001010100000;
   assign mem[141951:141920] = 32'b00000001000000000111011101110100;
   assign mem[141983:141952] = 32'b00000010100000000101110010010000;
   assign mem[142015:141984] = 32'b00000101111110110011000101100000;
   assign mem[142047:142016] = 32'b11110110110001110000011101100000;
   assign mem[142079:142048] = 32'b11111010001111100011000011001000;
   assign mem[142111:142080] = 32'b11111101010000100100000110010000;
   assign mem[142143:142112] = 32'b11111010110101010110101010111000;
   assign mem[142175:142144] = 32'b11111110100100100101011101011000;
   assign mem[142207:142176] = 32'b00000011110000011001101001001000;
   assign mem[142239:142208] = 32'b11111111101110000001110010000010;
   assign mem[142271:142240] = 32'b11111101011010010000110000010100;
   assign mem[142303:142272] = 32'b11111101000001000101001000000100;
   assign mem[142335:142304] = 32'b11111011101010000011010001110000;
   assign mem[142367:142336] = 32'b11111101010011010011110101100000;
   assign mem[142399:142368] = 32'b00000001100111100110001111011000;
   assign mem[142431:142400] = 32'b00000011110000100010000001111100;
   assign mem[142463:142432] = 32'b11111000111011111000000100110000;
   assign mem[142495:142464] = 32'b11111011101001110000100111011000;
   assign mem[142527:142496] = 32'b11110111100110010100001101000000;
   assign mem[142559:142528] = 32'b00000000101010111110110000010010;
   assign mem[142591:142560] = 32'b00000000101001010000001101011010;
   assign mem[142623:142592] = 32'b00000000111000000101010110100011;
   assign mem[142655:142624] = 32'b11111101010100111111000111100000;
   assign mem[142687:142656] = 32'b00000010011000011011010001100100;
   assign mem[142719:142688] = 32'b00000100111111010110100010010000;
   assign mem[142751:142720] = 32'b00000001000001110011001101011000;
   assign mem[142783:142752] = 32'b00000000001110100001011100010010;
   assign mem[142815:142784] = 32'b00000000010010100000101100010100;
   assign mem[142847:142816] = 32'b11110110011101101001101011100000;
   assign mem[142879:142848] = 32'b00000110001101111001110001101000;
   assign mem[142911:142880] = 32'b00000110001110111001001111111000;
   assign mem[142943:142912] = 32'b00000010000100110011000111100000;
   assign mem[142975:142944] = 32'b00000011010110011000100010001100;
   assign mem[143007:142976] = 32'b00000011000001000000110111010100;
   assign mem[143039:143008] = 32'b11111110101100010001001011011010;
   assign mem[143071:143040] = 32'b00000100110100010010011001001000;
   assign mem[143103:143072] = 32'b11111010011010111001110110011000;
   assign mem[143135:143104] = 32'b11111100110100110101000101000100;
   assign mem[143167:143136] = 32'b11110010100100111000011100110000;
   assign mem[143199:143168] = 32'b00000011010110111111011100111000;
   assign mem[143231:143200] = 32'b00000100010110110001110001011000;
   assign mem[143263:143232] = 32'b00000011001100010111001100001100;
   assign mem[143295:143264] = 32'b00001001010011010111000001000000;
   assign mem[143327:143296] = 32'b00000001011100001110101111001110;
   assign mem[143359:143328] = 32'b00000011101111110001011101111100;
   assign mem[143391:143360] = 32'b11111010001110101101111101011000;
   assign mem[143423:143392] = 32'b11101101111111001101000010000000;
   assign mem[143455:143424] = 32'b11111111101010000110111001000101;
   assign mem[143487:143456] = 32'b11111101101010011001010001111000;
   assign mem[143519:143488] = 32'b00000011001110010111010011100100;
   assign mem[143551:143520] = 32'b11111110001100000101101111111000;
   assign mem[143583:143552] = 32'b00000100100111011110101011000000;
   assign mem[143615:143584] = 32'b11111101010001111001110001010000;
   assign mem[143647:143616] = 32'b00000011101100110111001111110000;
   assign mem[143679:143648] = 32'b00000100011010001111001010110000;
   assign mem[143711:143680] = 32'b11111101000010010110111110000100;
   assign mem[143743:143712] = 32'b00001100011011111000000111000000;
   assign mem[143775:143744] = 32'b00000111010100101001010011001000;
   assign mem[143807:143776] = 32'b11111000001001111110010110011000;
   assign mem[143839:143808] = 32'b00000110010111011010111011010000;
   assign mem[143871:143840] = 32'b11111110110110011001000100111110;
   assign mem[143903:143872] = 32'b11111001000110001010100100111000;
   assign mem[143935:143904] = 32'b00000000001101011010000011011011;
   assign mem[143967:143936] = 32'b11101011111101011000111100100000;
   assign mem[143999:143968] = 32'b11100011100101010101110010100000;
   assign mem[144031:144000] = 32'b00000101110011000111101000111000;
   assign mem[144063:144032] = 32'b00000000110101010111111010000010;
   assign mem[144095:144064] = 32'b00000001000001111010101100100010;
   assign mem[144127:144096] = 32'b11111101011111111100000001010000;
   assign mem[144159:144128] = 32'b11110011000110000000110110100000;
   assign mem[144191:144160] = 32'b11111100110011101111001000101000;
   assign mem[144223:144192] = 32'b11111111011110011110101011110011;
   assign mem[144255:144224] = 32'b11111011011010011010101010110000;
   assign mem[144287:144256] = 32'b00001001000011000010001111000000;
   assign mem[144319:144288] = 32'b00000101111010010100101110101000;
   assign mem[144351:144320] = 32'b11111001000111011101111010110000;
   assign mem[144383:144352] = 32'b00000011111010010110010100101000;
   assign mem[144415:144384] = 32'b00000100010001111010100000110000;
   assign mem[144447:144416] = 32'b00000111000100010100101111101000;
   assign mem[144479:144448] = 32'b11111100000111000000100011100100;
   assign mem[144511:144480] = 32'b11111101101101011010101011100100;
   assign mem[144543:144512] = 32'b11110110000110010000011101100000;
   assign mem[144575:144544] = 32'b00001001010001100010000110000000;
   assign mem[144607:144576] = 32'b11111011100011001011101001111000;
   assign mem[144639:144608] = 32'b11111110100100101101110000001110;
   assign mem[144671:144640] = 32'b11111100010100101101011111011100;
   assign mem[144703:144672] = 32'b00000000111010001000100001010101;
   assign mem[144735:144704] = 32'b00000111100111111101000010000000;
   assign mem[144767:144736] = 32'b11111111101100001110110011111001;
   assign mem[144799:144768] = 32'b11110100011011111110000001010000;
   assign mem[144831:144800] = 32'b11111100101000111010011101101000;
   assign mem[144863:144832] = 32'b11111100101111001000100100100100;
   assign mem[144895:144864] = 32'b00000111111011110110001100000000;
   assign mem[144927:144896] = 32'b11110011101110101100000111110000;
   assign mem[144959:144928] = 32'b00000000011011010111101000011101;
   assign mem[144991:144960] = 32'b00000010111110000011010000111100;
   assign mem[145023:144992] = 32'b11111011000110101011110111001000;
   assign mem[145055:145024] = 32'b11111010111101111000001110100000;
   assign mem[145087:145056] = 32'b11111011010110101111111001110000;
   assign mem[145119:145088] = 32'b00000011010100011100110011010100;
   assign mem[145151:145120] = 32'b11111100110000110110110000111100;
   assign mem[145183:145152] = 32'b00000001110100011000111100000110;
   assign mem[145215:145184] = 32'b11111010001010001100011100101000;
   assign mem[145247:145216] = 32'b00000100010101000110101110001000;
   assign mem[145279:145248] = 32'b00000101011011100011111010010000;
   assign mem[145311:145280] = 32'b00000001011100101101111100001000;
   assign mem[145343:145312] = 32'b11111110101000010011011001001110;
   assign mem[145375:145344] = 32'b11111100000100011100001000001100;
   assign mem[145407:145376] = 32'b11111001011011101001100000110000;
   assign mem[145439:145408] = 32'b00000111011010111010111110110000;
   assign mem[145471:145440] = 32'b00000011011001000001000100100100;
   assign mem[145503:145472] = 32'b00001001001010101101010110010000;
   assign mem[145535:145504] = 32'b11111110110111011111000110000100;
   assign mem[145567:145536] = 32'b11111101011110000010000100000100;
   assign mem[145599:145568] = 32'b11110110110110111001010101100000;
   assign mem[145631:145600] = 32'b00000011000001000111111101100100;
   assign mem[145663:145632] = 32'b11111111010111010001001110000011;
   assign mem[145695:145664] = 32'b00001000100101110111001100000000;
   assign mem[145727:145696] = 32'b11111100010101100011000101010000;
   assign mem[145759:145728] = 32'b00000010100111110000010011110100;
   assign mem[145791:145760] = 32'b11111010111110010100001000001000;
   assign mem[145823:145792] = 32'b00000101001000011010111100010000;
   assign mem[145855:145824] = 32'b11111111010100000000011001101100;
   assign mem[145887:145856] = 32'b00000000000111110010110101100011;
   assign mem[145919:145888] = 32'b00000010111010001010010101100100;
   assign mem[145951:145920] = 32'b00000110110001111101100110000000;
   assign mem[145983:145952] = 32'b11111000011101010110011010000000;
   assign mem[146015:145984] = 32'b00001000010001010100101101110000;
   assign mem[146047:146016] = 32'b11111111110110001000001110111011;
   assign mem[146079:146048] = 32'b11111000000001000100111001001000;
   assign mem[146111:146080] = 32'b11111001000010001111100010011000;
   assign mem[146143:146112] = 32'b11111000100101101000110011010000;
   assign mem[146175:146144] = 32'b00000110000111000100110111110000;
   assign mem[146207:146176] = 32'b11111110111010110010011000001110;
   assign mem[146239:146208] = 32'b11111110101110011110010110100010;
   assign mem[146271:146240] = 32'b11110111111111011100100100100000;
   assign mem[146303:146272] = 32'b00000011010110101011000101000100;
   assign mem[146335:146304] = 32'b00000011010001111011000000010000;
   assign mem[146367:146336] = 32'b11110011110011010100101111000000;
   assign mem[146399:146368] = 32'b11111101111111000001100000100100;
   assign mem[146431:146400] = 32'b00000110100010011101111110011000;
   assign mem[146463:146432] = 32'b00000010110000101011001101000000;
   assign mem[146495:146464] = 32'b11111111111000001001111111010101;
   assign mem[146527:146496] = 32'b11111111010011111010000000001110;
   assign mem[146559:146528] = 32'b00000010110111110100111111010000;
   assign mem[146591:146560] = 32'b11111100000100001111001001011100;
   assign mem[146623:146592] = 32'b00000001100010010100001000011000;
   assign mem[146655:146624] = 32'b11111101011100100011000011101000;
   assign mem[146687:146656] = 32'b00000001111100110001001101010110;
   assign mem[146719:146688] = 32'b11111111101011000100010110101100;
   assign mem[146751:146720] = 32'b11111011010111111100101001001000;
   assign mem[146783:146752] = 32'b11111010111011001110111100010000;
   assign mem[146815:146784] = 32'b00000010101001111000001101001100;
   assign mem[146847:146816] = 32'b11111111111011000011000111001100;
   assign mem[146879:146848] = 32'b00000000101111101001001100100100;
   assign mem[146911:146880] = 32'b00000100110000100001000010101000;
   assign mem[146943:146912] = 32'b11111101000101000001111101101100;
   assign mem[146975:146944] = 32'b00000010011101000001100001110100;
   assign mem[147007:146976] = 32'b11111100111000100111100010100100;
   assign mem[147039:147008] = 32'b11110011000100100001100111100000;
   assign mem[147071:147040] = 32'b00000011010000001110110000111000;
   assign mem[147103:147072] = 32'b11110000100010010011110010010000;
   assign mem[147135:147104] = 32'b00000100111011111100001111101000;
   assign mem[147167:147136] = 32'b00001001001100101001010001010000;
   assign mem[147199:147168] = 32'b00001000101110001001010110100000;
   assign mem[147231:147200] = 32'b11111000101001010100000011101000;
   assign mem[147263:147232] = 32'b11110000100110000111001101000000;
   assign mem[147295:147264] = 32'b00000010001111110001010010101100;
   assign mem[147327:147296] = 32'b11111111010010101010100111010111;
   assign mem[147359:147328] = 32'b00000110001110110001011110111000;
   assign mem[147391:147360] = 32'b11111110111110001011010101000000;
   assign mem[147423:147392] = 32'b00001001111101000011011000010000;
   assign mem[147455:147424] = 32'b00000110101001011111100011011000;
   assign mem[147487:147456] = 32'b00000100101000011000011101001000;
   assign mem[147519:147488] = 32'b11111010001110010110000111001000;
   assign mem[147551:147520] = 32'b00000111001010111010111001001000;
   assign mem[147583:147552] = 32'b00000101000100111100111110010000;
   assign mem[147615:147584] = 32'b00001000111001010100101010110000;
   assign mem[147647:147616] = 32'b11111011010011011001001010001000;
   assign mem[147679:147648] = 32'b11111100000100111001001111110000;
   assign mem[147711:147680] = 32'b11111111111100000111111010110011;
   assign mem[147743:147712] = 32'b00000000111101110001010000111000;
   assign mem[147775:147744] = 32'b00000011110111111000111111000100;
   assign mem[147807:147776] = 32'b00000001111000110110100000110010;
   assign mem[147839:147808] = 32'b11110110011100111011111011110000;
   assign mem[147871:147840] = 32'b11111011101101010110111100110000;
   assign mem[147903:147872] = 32'b11111010011010100110011100001000;
   assign mem[147935:147904] = 32'b11111011111011111111111010000000;
   assign mem[147967:147936] = 32'b11111010001000010110100100110000;
   assign mem[147999:147968] = 32'b11111110100010010100011111101100;
   assign mem[148031:148000] = 32'b11111111100011001011110111010010;
   assign mem[148063:148032] = 32'b11111110010101000101100010100000;
   assign mem[148095:148064] = 32'b11110110111010111110111110000000;
   assign mem[148127:148096] = 32'b00000100011110100110100110111000;
   assign mem[148159:148128] = 32'b00000111111111001001110101000000;
   assign mem[148191:148160] = 32'b11111101100101110111011001111100;
   assign mem[148223:148192] = 32'b00000011001010101010010110100000;
   assign mem[148255:148224] = 32'b11111111001011000011101111111011;
   assign mem[148287:148256] = 32'b00000000001101111100110110111100;
   assign mem[148319:148288] = 32'b11111110111000011001110101010100;
   assign mem[148351:148320] = 32'b11111101000110011110101100110000;
   assign mem[148383:148352] = 32'b00001000100111011001110011010000;
   assign mem[148415:148384] = 32'b11111110001011100011101001001010;
   assign mem[148447:148416] = 32'b11111100011010010100011000001100;
   assign mem[148479:148448] = 32'b11111111111000110000100010110110;
   assign mem[148511:148480] = 32'b11111110111000111001111100011110;
   assign mem[148543:148512] = 32'b11111100111100011101001000110100;
   assign mem[148575:148544] = 32'b00001000010011111011101001010000;
   assign mem[148607:148576] = 32'b11111111100111110101011011000010;
   assign mem[148639:148608] = 32'b11111010100001001111110111011000;
   assign mem[148671:148640] = 32'b00000100011000000000100110101000;
   assign mem[148703:148672] = 32'b11111001110010101010011101110000;
   assign mem[148735:148704] = 32'b00000100110100110001011100001000;
   assign mem[148767:148736] = 32'b11111101100110001110011101100100;
   assign mem[148799:148768] = 32'b11111100100111101101111100000000;
   assign mem[148831:148800] = 32'b00000001010011000110100001010100;
   assign mem[148863:148832] = 32'b00000010010010100101001111010000;
   assign mem[148895:148864] = 32'b11111101101101100010011011010000;
   assign mem[148927:148896] = 32'b00000010111000011110111101111100;
   assign mem[148959:148928] = 32'b11110100000111001000000010010000;
   assign mem[148991:148960] = 32'b11111110100001001111110110010110;
   assign mem[149023:148992] = 32'b11101100010100101110100010100000;
   assign mem[149055:149024] = 32'b00000011110011101100001100000000;
   assign mem[149087:149056] = 32'b00000101010111011100000110110000;
   assign mem[149119:149088] = 32'b00000010101010101101100010101000;
   assign mem[149151:149120] = 32'b11111110100110111111011101001000;
   assign mem[149183:149152] = 32'b00010111010011000101000000100000;
   assign mem[149215:149184] = 32'b00000100000100011001100001000000;
   assign mem[149247:149216] = 32'b11110001000000101000011001110000;
   assign mem[149279:149248] = 32'b11110000000000011001010001000000;
   assign mem[149311:149280] = 32'b00001101000110010010001111000000;
   assign mem[149343:149312] = 32'b11111100110111101100001010101000;
   assign mem[149375:149344] = 32'b00000101100010000011101110011000;
   assign mem[149407:149376] = 32'b00000010011001101010110111010100;
   assign mem[149439:149408] = 32'b00000001000111100011001011000010;
   assign mem[149471:149440] = 32'b11111110010001000010011001011010;
   assign mem[149503:149472] = 32'b00000011000000011101101101010100;
   assign mem[149535:149504] = 32'b11111011100101110000100110100000;
   assign mem[149567:149536] = 32'b00000101101101011111011001101000;
   assign mem[149599:149568] = 32'b11111111100010010110001010101011;
   assign mem[149631:149600] = 32'b11111110101010000001101011111000;
   assign mem[149663:149632] = 32'b11111100011011000011010011111100;
   assign mem[149695:149664] = 32'b11110110100010110000111000100000;
   assign mem[149727:149696] = 32'b00000010001111000010111010011000;
   assign mem[149759:149728] = 32'b00000011010011000001000111100000;
   assign mem[149791:149760] = 32'b11111010110001100110110010110000;
   assign mem[149823:149792] = 32'b00000000100000011110111010010100;
   assign mem[149855:149824] = 32'b11111100101101010111010100010100;
   assign mem[149887:149856] = 32'b11110111101001100000100111000000;
   assign mem[149919:149888] = 32'b00000001101100000010010000111110;
   assign mem[149951:149920] = 32'b00000101111101101010010010000000;
   assign mem[149983:149952] = 32'b11111101010110010010010011011000;
   assign mem[150015:149984] = 32'b00000101010011000101100100110000;
   assign mem[150047:150016] = 32'b00000000001000011100010010110101;
   assign mem[150079:150048] = 32'b11111110011111001001010110110110;
   assign mem[150111:150080] = 32'b11111001010000000001000101011000;
   assign mem[150143:150112] = 32'b00000100100111000100001001100000;
   assign mem[150175:150144] = 32'b11111010011101101010110011101000;
   assign mem[150207:150176] = 32'b00000000111000011101000011111110;
   assign mem[150239:150208] = 32'b00000000010100101001100111110100;
   assign mem[150271:150240] = 32'b00000001110111110110101100011100;
   assign mem[150303:150272] = 32'b00000001001110000001110111001110;
   assign mem[150335:150304] = 32'b00000000001110011000111110011101;
   assign mem[150367:150336] = 32'b11111101101000010111001110111000;
   assign mem[150399:150368] = 32'b11111111101111110010000110000010;
   assign mem[150431:150400] = 32'b00000001011011111110101011001010;
   assign mem[150463:150432] = 32'b11111111011101010011011001011010;
   assign mem[150495:150464] = 32'b11111110011010101111010010001100;
   assign mem[150527:150496] = 32'b00000010101101110010000011101100;
   assign mem[150559:150528] = 32'b00000010100001000011111001110000;
   assign mem[150591:150560] = 32'b11111011101101011000000110111000;
   assign mem[150623:150592] = 32'b00000000000110010011100110001000;
   assign mem[150655:150624] = 32'b11111000110000011111011001010000;
   assign mem[150687:150656] = 32'b11111111100111001001101110111011;
   assign mem[150719:150688] = 32'b00000011000001001001011000000100;
   assign mem[150751:150720] = 32'b11111110000000010100000110111010;
   assign mem[150783:150752] = 32'b00000010100111011101010011000100;
   assign mem[150815:150784] = 32'b00000001111100000010000100110110;
   assign mem[150847:150816] = 32'b11111001100101111110011001100000;
   assign mem[150879:150848] = 32'b11111110001111001010010010110100;
   assign mem[150911:150880] = 32'b00000000111101101000001011111011;
   assign mem[150943:150912] = 32'b11101011110011001101100110000000;
   assign mem[150975:150944] = 32'b11111011100011011000100100110000;
   assign mem[151007:150976] = 32'b00001100101100100101010110100000;
   assign mem[151039:151008] = 32'b00000101100010100000000010011000;
   assign mem[151071:151040] = 32'b11111011100111000011101000100000;
   assign mem[151103:151072] = 32'b11111110110010101011101011110110;
   assign mem[151135:151104] = 32'b11111101010010010111100110110100;
   assign mem[151167:151136] = 32'b11110110100010001111110000100000;
   assign mem[151199:151168] = 32'b00000011100000111101111110110000;
   assign mem[151231:151200] = 32'b11111111110011000111001011101101;
   assign mem[151263:151232] = 32'b11101101001101001111100100000000;
   assign mem[151295:151264] = 32'b11111001101011000001010111110000;
   assign mem[151327:151296] = 32'b00001001111011011010111010010000;
   assign mem[151359:151328] = 32'b00000101010010001100110100101000;
   assign mem[151391:151360] = 32'b11111111110110000010010010001000;
   assign mem[151423:151392] = 32'b00001011111101011011100110010000;
   assign mem[151455:151424] = 32'b00000000111111110100010011000100;
   assign mem[151487:151456] = 32'b11111101011000001000101101010000;
   assign mem[151519:151488] = 32'b00000110100101111010011010010000;
   assign mem[151551:151520] = 32'b00000001010110110001101100001100;
   assign mem[151583:151552] = 32'b00000101110111001011111000010000;
   assign mem[151615:151584] = 32'b11111111010111110101010110111101;
   assign mem[151647:151616] = 32'b11110111001010100000101010000000;
   assign mem[151679:151648] = 32'b11111011011001000110001011100000;
   assign mem[151711:151680] = 32'b00000000001011101001111101101000;
   assign mem[151743:151712] = 32'b11110110111000101011001000100000;
   assign mem[151775:151744] = 32'b00000101000100101110010100001000;
   assign mem[151807:151776] = 32'b11101101110100101000011011100000;
   assign mem[151839:151808] = 32'b00000110110001010111110011101000;
   assign mem[151871:151840] = 32'b00000000000001111000110011001110;
   assign mem[151903:151872] = 32'b00000010101000010001000111110100;
   assign mem[151935:151904] = 32'b11111111001110111011110000101010;
   assign mem[151967:151936] = 32'b11111110001110111001100110010000;
   assign mem[151999:151968] = 32'b11111110000010111100010101100110;
   assign mem[152031:152000] = 32'b00000110100001010001101101010000;
   assign mem[152063:152032] = 32'b00000011101100011011110011011100;
   assign mem[152095:152064] = 32'b11111101101010100011111111100000;
   assign mem[152127:152096] = 32'b11101111100011110110001110100000;
   assign mem[152159:152128] = 32'b11111101110000010010010101010000;
   assign mem[152191:152160] = 32'b00001000010000111001000010010000;
   assign mem[152223:152192] = 32'b00001001010001010101000110100000;
   assign mem[152255:152224] = 32'b11111100010001010101011001011000;
   assign mem[152287:152256] = 32'b11110111001110001100100000100000;
   assign mem[152319:152288] = 32'b11111111101001001101000001010100;
   assign mem[152351:152320] = 32'b11111110001100101011110111101000;
   assign mem[152383:152352] = 32'b11111100111101100011101001111000;
   assign mem[152415:152384] = 32'b11111100110111111011100010001000;
   assign mem[152447:152416] = 32'b00000101101011010001011010011000;
   assign mem[152479:152448] = 32'b00000001101010010000011010101110;
   assign mem[152511:152480] = 32'b11111110010000011000001010011110;
   assign mem[152543:152512] = 32'b11111101110101100110110010110100;
   assign mem[152575:152544] = 32'b11111110000110001001111100011010;
   assign mem[152607:152576] = 32'b00000000100101101111100011000110;
   assign mem[152639:152608] = 32'b00001010000000111110011010100000;
   assign mem[152671:152640] = 32'b00000110110100110011011110100000;
   assign mem[152703:152672] = 32'b11111000000000110100110100101000;
   assign mem[152735:152704] = 32'b00000011001101100001100000110100;
   assign mem[152767:152736] = 32'b00000000010100110000100111001001;
   assign mem[152799:152768] = 32'b11110101001001101001000100000000;
   assign mem[152831:152800] = 32'b11111110000000000011110011001000;
   assign mem[152863:152832] = 32'b11101110010011001011011000100000;
   assign mem[152895:152864] = 32'b00001010001100100100000010110000;
   assign mem[152927:152896] = 32'b00000010001100111110011001110100;
   assign mem[152959:152928] = 32'b00000110000101000101000010001000;
   assign mem[152991:152960] = 32'b11111011010001010001000100010000;
   assign mem[153023:152992] = 32'b00000011010101010001101011000000;
   assign mem[153055:153024] = 32'b11111111100011111001001001011100;
   assign mem[153087:153056] = 32'b11110110111000001010110000100000;
   assign mem[153119:153088] = 32'b00000010111100010100110101111100;
   assign mem[153151:153120] = 32'b00000011011111010001110110011100;
   assign mem[153183:153152] = 32'b00000100010111011101100010111000;
   assign mem[153215:153184] = 32'b00000010001010111101000100101100;
   assign mem[153247:153216] = 32'b11110111011101001001110110010000;
   assign mem[153279:153248] = 32'b11111000110010000100000010111000;
   assign mem[153311:153280] = 32'b11111100011011111011001000111100;
   assign mem[153343:153312] = 32'b00000011011001000000000110100100;
   assign mem[153375:153344] = 32'b00000100011111100010010010111000;
   assign mem[153407:153376] = 32'b11111111011100001110000011000011;
   assign mem[153439:153408] = 32'b11111001001000010010010110100000;
   assign mem[153471:153440] = 32'b00000100011011011010110111111000;
   assign mem[153503:153472] = 32'b11110111001011011100000101010000;
   assign mem[153535:153504] = 32'b00000011100100010101101010011000;
   assign mem[153567:153536] = 32'b11111101010010000000111011010000;
   assign mem[153599:153568] = 32'b11111011101011111110010110010000;
   assign mem[153631:153600] = 32'b00000000110011001101000101101010;
   assign mem[153663:153632] = 32'b00000000011001001011000101101100;
   assign mem[153695:153664] = 32'b11111111001111011101110100001100;
   assign mem[153727:153696] = 32'b11111011100110001110010011101000;
   assign mem[153759:153728] = 32'b00000010011001110010011111101000;
   assign mem[153791:153760] = 32'b11111111010010001111000101110010;
   assign mem[153823:153792] = 32'b11111111011110101111100111011110;
   assign mem[153855:153824] = 32'b11111110001110111000111001001010;
   assign mem[153887:153856] = 32'b11111101111111011111010101111000;
   assign mem[153919:153888] = 32'b00000000111010110100101011111100;
   assign mem[153951:153920] = 32'b00000001001010010010001010111110;
   assign mem[153983:153952] = 32'b11111101010111110011111000011100;
   assign mem[154015:153984] = 32'b11111101000000011100110111101000;
   assign mem[154047:154016] = 32'b11110001011010010010101100000000;
   assign mem[154079:154048] = 32'b00000000001110111010011010100110;
   assign mem[154111:154080] = 32'b00000101001101101001110101010000;
   assign mem[154143:154112] = 32'b00000011110101000001000010100100;
   assign mem[154175:154144] = 32'b11111101011100010001010011000000;
   assign mem[154207:154176] = 32'b11111011011101011010100110001000;
   assign mem[154239:154208] = 32'b00000000011100000101000110001010;
   assign mem[154271:154240] = 32'b00000011000000110011100101111000;
   assign mem[154303:154272] = 32'b11110110010100111111011111010000;
   assign mem[154335:154304] = 32'b00000010010010101111100101011000;
   assign mem[154367:154336] = 32'b11111100111101011001011010110000;
   assign mem[154399:154368] = 32'b11110100001101011110100011000000;
   assign mem[154431:154400] = 32'b00000010110001101011111010001000;
   assign mem[154463:154432] = 32'b11111100000100101101011100111000;
   assign mem[154495:154464] = 32'b00000110101100111101010100000000;
   assign mem[154527:154496] = 32'b00000000010100111000111110010001;
   assign mem[154559:154528] = 32'b00000000010011101110101000001010;
   assign mem[154591:154560] = 32'b00000010011100011101101101101000;
   assign mem[154623:154592] = 32'b00001100101110011111111010100000;
   assign mem[154655:154624] = 32'b00001001000001010001110010000000;
   assign mem[154687:154656] = 32'b11111101000010001011000110011000;
   assign mem[154719:154688] = 32'b00000101001101010001011010101000;
   assign mem[154751:154720] = 32'b00000000010011110001000101110011;
   assign mem[154783:154752] = 32'b00001000010010100101011000100000;
   assign mem[154815:154784] = 32'b11101000100000011000010100000000;
   assign mem[154847:154816] = 32'b11110111110100100111110111010000;
   assign mem[154879:154848] = 32'b11111010010110010100000100010000;
   assign mem[154911:154880] = 32'b11111110110001010100001010110110;
   assign mem[154943:154912] = 32'b11111011000111010110000101110000;
   assign mem[154975:154944] = 32'b00000010110111010110110100111000;
   assign mem[155007:154976] = 32'b11111001101000011100101100011000;
   assign mem[155039:155008] = 32'b11111001101101001111001000101000;
   assign mem[155071:155040] = 32'b00000101100000110011111100000000;
   assign mem[155103:155072] = 32'b00000010010010011000111111101000;
   assign mem[155135:155104] = 32'b00000011101001101000001100110000;
   assign mem[155167:155136] = 32'b00000010110011101110100011001000;
   assign mem[155199:155168] = 32'b11110100001110100001111000100000;
   assign mem[155231:155200] = 32'b00000010010110111110110110011000;
   assign mem[155263:155232] = 32'b11111000111000011011000011101000;
   assign mem[155295:155264] = 32'b11111111000000111110000011101111;
   assign mem[155327:155296] = 32'b11111110000000111110100110100100;
   assign mem[155359:155328] = 32'b11110110100010101011101010100000;
   assign mem[155391:155360] = 32'b11111110000010010101110100010100;
   assign mem[155423:155392] = 32'b11110110100010011111110100000000;
   assign mem[155455:155424] = 32'b00000011010001111001111111011100;
   assign mem[155487:155456] = 32'b00000101111000110111111111111000;
   assign mem[155519:155488] = 32'b00001001011100000111101011000000;
   assign mem[155551:155520] = 32'b11111110011111110101111101101110;
   assign mem[155583:155552] = 32'b00000100000000000001110110011000;
   assign mem[155615:155584] = 32'b11111111000101011111111111001000;
   assign mem[155647:155616] = 32'b11111001001100111001111110100000;
   assign mem[155679:155648] = 32'b00000011011000101001010100110100;
   assign mem[155711:155680] = 32'b00000111000000101100111110100000;
   assign mem[155743:155712] = 32'b11111101111111000110010101111100;
   assign mem[155775:155744] = 32'b00000100010111110001000001001000;
   assign mem[155807:155776] = 32'b11111100101110100100000011000100;
   assign mem[155839:155808] = 32'b00000101010001010011010001011000;
   assign mem[155871:155840] = 32'b11111011100001001110100100111000;
   assign mem[155903:155872] = 32'b00000101101000010000101011100000;
   assign mem[155935:155904] = 32'b00000000110010111100110111110000;
   assign mem[155967:155936] = 32'b00001001000111110110000001010000;
   assign mem[155999:155968] = 32'b11110101010110011010001000100000;
   assign mem[156031:156000] = 32'b11111000011111001001000110001000;
   assign mem[156063:156032] = 32'b11111010001011000101111011010000;
   assign mem[156095:156064] = 32'b00001000111010010011101110000000;
   assign mem[156127:156096] = 32'b11101110011100111000001000000000;
   assign mem[156159:156128] = 32'b11110101001110100111000010100000;
   assign mem[156191:156160] = 32'b00000110001100111101110000100000;
   assign mem[156223:156192] = 32'b11111100011101110100111101100000;
   assign mem[156255:156224] = 32'b00000101110010001101100110001000;
   assign mem[156287:156256] = 32'b11111000011111110001110100110000;
   assign mem[156319:156288] = 32'b11110000011110011101001111000000;
   assign mem[156351:156320] = 32'b00000001100100000000011000101010;
   assign mem[156383:156352] = 32'b11111001010111111100011101011000;
   assign mem[156415:156384] = 32'b00000100011110010111110110010000;
   assign mem[156447:156416] = 32'b00001000110100001011001100000000;
   assign mem[156479:156448] = 32'b00000001011111011111111000000000;
   assign mem[156511:156480] = 32'b11110110001111001110111000110000;
   assign mem[156543:156512] = 32'b11111110011101110000010110000100;
   assign mem[156575:156544] = 32'b00000010111010111101110101011100;
   assign mem[156607:156576] = 32'b00000000001011101101101001101100;
   assign mem[156639:156608] = 32'b11111110111011000011010101001000;
   assign mem[156671:156640] = 32'b00000011000010010111101100001100;
   assign mem[156703:156672] = 32'b00000011100111000010101010001100;
   assign mem[156735:156704] = 32'b00000110110010111001100100100000;
   assign mem[156767:156736] = 32'b11111100101011100010010100110000;
   assign mem[156799:156768] = 32'b11111100010010110110100011001000;
   assign mem[156831:156800] = 32'b11111111100010100110010110000101;
   assign mem[156863:156832] = 32'b00000100000100000100101001110000;
   assign mem[156895:156864] = 32'b00000100100000000101010111110000;
   assign mem[156927:156896] = 32'b00000011111110111011110111010000;
   assign mem[156959:156928] = 32'b11110000011111111101001000000000;
   assign mem[156991:156960] = 32'b11110111010100001000000011110000;
   assign mem[157023:156992] = 32'b11111101111010101101110101110000;
   assign mem[157055:157024] = 32'b00000110100001010100111001110000;
   assign mem[157087:157056] = 32'b11110011101000001010111101010000;
   assign mem[157119:157088] = 32'b11111001101100110000111111001000;
   assign mem[157151:157120] = 32'b11110110110100100011110100110000;
   assign mem[157183:157152] = 32'b00000001110000100111011010011010;
   assign mem[157215:157184] = 32'b00000110100000101000111000001000;
   assign mem[157247:157216] = 32'b00000010110010110101010100000000;
   assign mem[157279:157248] = 32'b00001011100101101100011010000000;
   assign mem[157311:157280] = 32'b11111011001001001000101111011000;
   assign mem[157343:157312] = 32'b11111100000110001011010110001100;
   assign mem[157375:157344] = 32'b00000101100000100010101111010000;
   assign mem[157407:157376] = 32'b11110101000010111110111011100000;
   assign mem[157439:157408] = 32'b11110001111010011000000110000000;
   assign mem[157471:157440] = 32'b11111100010001010001000000010100;
   assign mem[157503:157472] = 32'b00000010000000011011111010010100;
   assign mem[157535:157504] = 32'b11111100101110100100111101110100;
   assign mem[157567:157536] = 32'b11111011000100100010100101000000;
   assign mem[157599:157568] = 32'b11111110000111101100110010010110;
   assign mem[157631:157600] = 32'b00001000001000111100111010010000;
   assign mem[157663:157632] = 32'b00000011001110001111101100001100;
   assign mem[157695:157664] = 32'b11110101100110011000011111110000;
   assign mem[157727:157696] = 32'b11111110010101110000110001111110;
   assign mem[157759:157728] = 32'b00000101010100001011101101000000;
   assign mem[157791:157760] = 32'b00000010011001111110110000111000;
   assign mem[157823:157792] = 32'b00000000010101101100010110101000;
   assign mem[157855:157824] = 32'b00000111000010000001011100001000;
   assign mem[157887:157856] = 32'b11111111000111010000110010111010;
   assign mem[157919:157888] = 32'b11110110110000001100011000010000;
   assign mem[157951:157920] = 32'b11111001110011010001011001101000;
   assign mem[157983:157952] = 32'b11111000100111101110011100110000;
   assign mem[158015:157984] = 32'b00000101100110100011010101100000;
   assign mem[158047:158016] = 32'b11111101010100000101001000110100;
   assign mem[158079:158048] = 32'b00000110001010111100100100010000;
   assign mem[158111:158080] = 32'b11110001110110011010001010010000;
   assign mem[158143:158112] = 32'b00000010110110010111100110010100;
   assign mem[158175:158144] = 32'b00000100000110111100001101011000;
   assign mem[158207:158176] = 32'b00000001011001011110001000001100;
   assign mem[158239:158208] = 32'b11111100001111100101100111001000;
   assign mem[158271:158240] = 32'b11110111011001011000111110110000;
   assign mem[158303:158272] = 32'b11111000001101010011100101110000;
   assign mem[158335:158304] = 32'b00000111101011010001010001011000;
   assign mem[158367:158336] = 32'b00000010111000101100001101110000;
   assign mem[158399:158368] = 32'b11111100011111111000010111010100;
   assign mem[158431:158400] = 32'b11111011101101000100110100001000;
   assign mem[158463:158432] = 32'b11111111000011111000000000111000;
   assign mem[158495:158464] = 32'b11111110111000000100011111101000;
   assign mem[158527:158496] = 32'b11111101101100111101110111111000;
   assign mem[158559:158528] = 32'b11111101011110101010101100100100;
   assign mem[158591:158560] = 32'b00000010001001001110111100111100;
   assign mem[158623:158592] = 32'b00000001010010111011010100101010;
   assign mem[158655:158624] = 32'b00000001100000100101001110010100;
   assign mem[158687:158656] = 32'b00000000100011000000101111110000;
   assign mem[158719:158688] = 32'b00000000010000100111101010110001;
   assign mem[158751:158720] = 32'b00000111000101111011100000101000;
   assign mem[158783:158752] = 32'b11111010010011101010011000101000;
   assign mem[158815:158784] = 32'b00000010111001010101000111100000;
   assign mem[158847:158816] = 32'b00000010001110101001001000001000;
   assign mem[158879:158848] = 32'b11110010110101100100001001100000;
   assign mem[158911:158880] = 32'b00000001110010110001110100001110;
   assign mem[158943:158912] = 32'b11111100111011001011111110101000;
   assign mem[158975:158944] = 32'b00000100000111001001000111100000;
   assign mem[159007:158976] = 32'b00000000010101111010000000100111;
   assign mem[159039:159008] = 32'b11111110000101101001011111010100;
   assign mem[159071:159040] = 32'b00000010100101001111001001111100;
   assign mem[159103:159072] = 32'b00000011001110001111010010000100;
   assign mem[159135:159104] = 32'b11111111110000111100010101010111;
   assign mem[159167:159136] = 32'b11110001011110111101011111100000;
   assign mem[159199:159168] = 32'b11111101101111101000010101100000;
   assign mem[159231:159200] = 32'b00000000101010000001111001100100;
   assign mem[159263:159232] = 32'b00000011110011010010110010110000;
   assign mem[159295:159264] = 32'b11111110010101101111110001010000;
   assign mem[159327:159296] = 32'b11111001010110000011010101000000;
   assign mem[159359:159328] = 32'b00000010010011110011011001111100;
   assign mem[159391:159360] = 32'b00000001001011000000101000011010;
   assign mem[159423:159392] = 32'b11111111000001100111100100111110;
   assign mem[159455:159424] = 32'b11111000011000001011101100111000;
   assign mem[159487:159456] = 32'b00000010001000011000011100101100;
   assign mem[159519:159488] = 32'b00000010000100000100111111010000;
   assign mem[159551:159520] = 32'b11111100000111111110011101111000;
   assign mem[159583:159552] = 32'b00001001001100111000010111100000;
   assign mem[159615:159584] = 32'b11111010001010101111011010000000;
   assign mem[159647:159616] = 32'b11111101000010011000010101101100;
   assign mem[159679:159648] = 32'b00000100010011101011111110011000;
   assign mem[159711:159680] = 32'b11110011111001110001110001100000;
   assign mem[159743:159712] = 32'b00000111101110001010111000101000;
   assign mem[159775:159744] = 32'b00000110011000011111111101100000;
   assign mem[159807:159776] = 32'b11111101111001011111011101010100;
   assign mem[159839:159808] = 32'b11111101111100001011011111110100;
   assign mem[159871:159840] = 32'b11111001011000110001111000101000;
   assign mem[159903:159872] = 32'b11111101010000011101001001111000;
   assign mem[159935:159904] = 32'b11111110101100100111110000100000;
   assign mem[159967:159936] = 32'b11111111011010110101010111001110;
   assign mem[159999:159968] = 32'b11110011001001100100110011100000;
   assign mem[160031:160000] = 32'b11111101000011100011101101110000;
   assign mem[160063:160032] = 32'b11111010011101000101100110110000;
   assign mem[160095:160064] = 32'b00000000111111000011100100001110;
   assign mem[160127:160096] = 32'b00000001101000110010110101001110;
   assign mem[160159:160128] = 32'b11110100101011000011100001110000;
   assign mem[160191:160160] = 32'b11111110010010010111101111001110;
   assign mem[160223:160192] = 32'b11111010101100100011001001010000;
   assign mem[160255:160224] = 32'b00000001101011111011110110111100;
   assign mem[160287:160256] = 32'b11111111000001001011010000110110;
   assign mem[160319:160288] = 32'b00000011011010011000111011111000;
   assign mem[160351:160320] = 32'b11111000001000010111111001101000;
   assign mem[160383:160352] = 32'b11110100000011101110110000100000;
   assign mem[160415:160384] = 32'b00000000110011000011000010101100;
   assign mem[160447:160416] = 32'b00000000100101001011011110011100;
   assign mem[160479:160448] = 32'b11110100101101110101010011010000;
   assign mem[160511:160480] = 32'b00000010101000101100010100111100;
   assign mem[160543:160512] = 32'b11111101111100000010010010011100;
   assign mem[160575:160544] = 32'b00000011001111010011111100110100;
   assign mem[160607:160576] = 32'b00000000001000100000101110011110;
   assign mem[160639:160608] = 32'b00000110110011111100011110001000;
   assign mem[160671:160640] = 32'b11111111000000110010000111001101;
   assign mem[160703:160672] = 32'b11111110110001001010111110100000;
   assign mem[160735:160704] = 32'b00000111000111011100110011110000;
   assign mem[160767:160736] = 32'b00000000011001000100100101110011;
   assign mem[160799:160768] = 32'b11111001011000000110101001000000;
   assign mem[160831:160800] = 32'b11111111101010001000110010011111;
   assign mem[160863:160832] = 32'b11111110001100011100101010010100;
   assign mem[160895:160864] = 32'b00000010011001000101010000000100;
   assign mem[160927:160896] = 32'b11111100011100111101111000000000;
   assign mem[160959:160928] = 32'b11111011111000011111100111100000;
   assign mem[160991:160960] = 32'b11111101110101010101001000011000;
   assign mem[161023:160992] = 32'b00000001010110110110011110101110;
   assign mem[161055:161024] = 32'b00000010110101100000100010001000;
   assign mem[161087:161056] = 32'b11111100011111011111010000001000;
   assign mem[161119:161088] = 32'b00000111111010100010101111010000;
   assign mem[161151:161120] = 32'b11111101001001000110111011100000;
   assign mem[161183:161152] = 32'b00000010100111010000010100011100;
   assign mem[161215:161184] = 32'b11111010010011110101101110111000;
   assign mem[161247:161216] = 32'b00000001110100011111011111101110;
   assign mem[161279:161248] = 32'b00000010101010000100110001010100;
   assign mem[161311:161280] = 32'b00000100011101101000011110110000;
   assign mem[161343:161312] = 32'b00000111011010111000100100001000;
   assign mem[161375:161344] = 32'b00000010100000000000010000110000;
   assign mem[161407:161376] = 32'b00000011000000110111001110111100;
   assign mem[161439:161408] = 32'b00001000101100001000000111000000;
   assign mem[161471:161440] = 32'b11111110001001100101010111011000;
   assign mem[161503:161472] = 32'b11111101101100000011000100110000;
   assign mem[161535:161504] = 32'b00000000100100100010101001001010;
   assign mem[161567:161536] = 32'b00000000000110100101110100111001;
   assign mem[161599:161568] = 32'b11110000111010111000001001100000;
   assign mem[161631:161600] = 32'b11111101100010011100000101010000;
   assign mem[161663:161632] = 32'b11111111101101111001101010110100;
   assign mem[161695:161664] = 32'b00000101111011101100011001010000;
   assign mem[161727:161696] = 32'b00000101011010010010111010110000;
   assign mem[161759:161728] = 32'b11110010111011001001101011000000;
   assign mem[161791:161760] = 32'b11111100111011001100100011010100;
   assign mem[161823:161792] = 32'b11110111010011001000111100000000;
   assign mem[161855:161824] = 32'b00000011100110100011101011111000;
   assign mem[161887:161856] = 32'b00000011100010001101100100110100;
   assign mem[161919:161888] = 32'b11111111011101011010111101010000;
   assign mem[161951:161920] = 32'b00000101100110110110100111110000;
   assign mem[161983:161952] = 32'b11111101001100111111111001101100;
   assign mem[162015:161984] = 32'b00000011100101100011010100011100;
   assign mem[162047:162016] = 32'b11111101000010111011000110010000;
   assign mem[162079:162048] = 32'b00000011000110011001111100101100;
   assign mem[162111:162080] = 32'b11111110100000001011111000001010;
   assign mem[162143:162112] = 32'b11111110101111100000011101110010;
   assign mem[162175:162144] = 32'b00000110001100100001111100010000;
   assign mem[162207:162176] = 32'b11110110000011101000011101110000;
   assign mem[162239:162208] = 32'b11110101000000101011101101010000;
   assign mem[162271:162240] = 32'b00000000000100100101001101010110;
   assign mem[162303:162272] = 32'b11111111101111100010100010011001;
   assign mem[162335:162304] = 32'b00000000010100000110111101011100;
   assign mem[162367:162336] = 32'b11111100011010001001111001001100;
   assign mem[162399:162368] = 32'b00000010010111101001001000001100;
   assign mem[162431:162400] = 32'b11111101001110010000001000010000;
   assign mem[162463:162432] = 32'b11111000000100010111011001011000;
   assign mem[162495:162464] = 32'b00000110011100110000101110111000;
   assign mem[162527:162496] = 32'b11111111100100100001100000111110;
   assign mem[162559:162528] = 32'b00000000000110010001111011010001;
   assign mem[162591:162560] = 32'b00000010101100011010101110100100;
   assign mem[162623:162592] = 32'b00000011000010100101110111011000;
   assign mem[162655:162624] = 32'b11111101010000010010110100111000;
   assign mem[162687:162656] = 32'b00000100011111011111100001001000;
   assign mem[162719:162688] = 32'b11111110010110010001000111111100;
   assign mem[162751:162720] = 32'b11111110000000111111010110101000;
   assign mem[162783:162752] = 32'b00000100001101011100010100110000;
   assign mem[162815:162784] = 32'b00000000111011000111000000101110;
   assign mem[162847:162816] = 32'b11111000111000001001001110100000;
   assign mem[162879:162848] = 32'b00000010000101101000101100110000;
   assign mem[162911:162880] = 32'b00000110111111101100011010010000;
   assign mem[162943:162912] = 32'b00000001100100000000110101010000;
   assign mem[162975:162944] = 32'b00000000001000101001100000001100;
   assign mem[163007:162976] = 32'b11101011010101001010010011000000;
   assign mem[163039:163008] = 32'b11111110110001001010000100010000;
   assign mem[163071:163040] = 32'b00000010100001100110011100011100;
   assign mem[163103:163072] = 32'b00000100111110111010001101110000;
   assign mem[163135:163104] = 32'b11111010100111010011010101100000;
   assign mem[163167:163136] = 32'b11111101011100001000100000110000;
   assign mem[163199:163168] = 32'b11111101010110100011111110011000;
   assign mem[163231:163200] = 32'b11111011011101001100000111110000;
   assign mem[163263:163232] = 32'b00000100101000001001100100101000;
   assign mem[163295:163264] = 32'b00000010100101010111101111010100;
   assign mem[163327:163296] = 32'b11110110011000100000010000010000;
   assign mem[163359:163328] = 32'b00000100000101110111011011000000;
   assign mem[163391:163360] = 32'b00001010101011110000011010010000;
   assign mem[163423:163392] = 32'b00000001000010001011011111110010;
   assign mem[163455:163424] = 32'b11110100110001000110110101100000;
   assign mem[163487:163456] = 32'b00000000110111001000110001001011;
   assign mem[163519:163488] = 32'b11110101010010000110000010110000;
   assign mem[163551:163520] = 32'b11110101000011100001101010110000;
   assign mem[163583:163552] = 32'b00000010110100000100111001010000;
   assign mem[163615:163584] = 32'b00000001010001111000110011111110;
   assign mem[163647:163616] = 32'b11110110100001011100001100000000;
   assign mem[163679:163648] = 32'b00000001000011110000100111111100;
   assign mem[163711:163680] = 32'b00000101111110000100000100110000;
   assign mem[163743:163712] = 32'b00000001000110110001011011100010;
   assign mem[163775:163744] = 32'b11111110000011010100010100110100;
   assign mem[163807:163776] = 32'b11111100001100011100000100011100;
   assign mem[163839:163808] = 32'b11111011111000100101011101101000;
   assign mem[163871:163840] = 32'b11111011111001101100010010010000;
   assign mem[163903:163872] = 32'b11110011010100011010001111100000;
   assign mem[163935:163904] = 32'b11111011110110001100010011110000;
   assign mem[163967:163936] = 32'b00000101111011010111000001100000;
   assign mem[163999:163968] = 32'b11110100000111111111110111010000;
   assign mem[164031:164000] = 32'b00000000011010010000000011110010;
   assign mem[164063:164032] = 32'b00000011101000110100111111110100;
   assign mem[164095:164064] = 32'b11110101011101011111111011100000;
   assign mem[164127:164096] = 32'b00000111000110110010010010100000;
   assign mem[164159:164128] = 32'b00000101001000100111001111000000;
   assign mem[164191:164160] = 32'b00000111011100101001001001011000;
   assign mem[164223:164192] = 32'b00000001111100011010110001100110;
   assign mem[164255:164224] = 32'b00000100010100000101010100110000;
   assign mem[164287:164256] = 32'b00000101100000010010010010011000;
   assign mem[164319:164288] = 32'b11111011111000100010111000000000;
   assign mem[164351:164320] = 32'b11101101010100001100001001000000;
   assign mem[164383:164352] = 32'b11110101101111101111111001110000;
   assign mem[164415:164384] = 32'b11111110101000010011110001111010;
   assign mem[164447:164416] = 32'b11111001111010111011001100001000;
   assign mem[164479:164448] = 32'b00000011000100101100001100111100;
   assign mem[164511:164480] = 32'b00000100001010101101010101000000;
   assign mem[164543:164512] = 32'b11111101011100101010001001101000;
   assign mem[164575:164544] = 32'b00000001011100110110101001010100;
   assign mem[164607:164576] = 32'b11111101110100111110110010101100;
   assign mem[164639:164608] = 32'b11110110000000100101111010010000;
   assign mem[164671:164640] = 32'b00000000110001000010001010010010;
   assign mem[164703:164672] = 32'b11111010101111001110010100010000;
   assign mem[164735:164704] = 32'b11111111110111010011111001010010;
   assign mem[164767:164736] = 32'b11111110111011011001101010101000;
   assign mem[164799:164768] = 32'b11111110010110000011001111101100;
   assign mem[164831:164800] = 32'b11111011010011111000000011001000;
   assign mem[164863:164832] = 32'b11110000101110000101110110110000;
   assign mem[164895:164864] = 32'b11111011111110000101000011100000;
   assign mem[164927:164896] = 32'b00000010011000010000010000110100;
   assign mem[164959:164928] = 32'b11110101001011000111100111100000;
   assign mem[164991:164960] = 32'b00000110101011011111000010000000;
   assign mem[165023:164992] = 32'b11111100010001011111010000110100;
   assign mem[165055:165024] = 32'b00000111000000000000010111001000;
   assign mem[165087:165056] = 32'b11111110101111010101001011010000;
   assign mem[165119:165088] = 32'b00000100000000010111010010100000;
   assign mem[165151:165120] = 32'b11111101110111011101001000110100;
   assign mem[165183:165152] = 32'b11111110010100001001011000001100;
   assign mem[165215:165184] = 32'b11111111001001111100100100101001;
   assign mem[165247:165216] = 32'b11110011010001110111100100000000;
   assign mem[165279:165248] = 32'b11111011101011111110010011111000;
   assign mem[165311:165280] = 32'b00001100110100011101100100010000;
   assign mem[165343:165312] = 32'b00000110110100100000010100110000;
   assign mem[165375:165344] = 32'b11111010010001111011010101010000;
   assign mem[165407:165376] = 32'b11111001110011101100111010100000;
   assign mem[165439:165408] = 32'b00000010110110011011110110110000;
   assign mem[165471:165440] = 32'b11111100010101110001010000110000;
   assign mem[165503:165472] = 32'b00000010000110011111001001011000;
   assign mem[165535:165504] = 32'b00000001100110001110111101000100;
   assign mem[165567:165536] = 32'b11111111100100010100011100010101;
   assign mem[165599:165568] = 32'b00000101000000111000010111100000;
   assign mem[165631:165600] = 32'b11111001110111101001111000111000;
   assign mem[165663:165632] = 32'b00000101000000010001110001010000;
   assign mem[165695:165664] = 32'b11111010000110011001011111010000;
   assign mem[165727:165696] = 32'b11111101101110011111111001111000;
   assign mem[165759:165728] = 32'b00000001011000001010100100001000;
   assign mem[165791:165760] = 32'b11110101101101011111110101000000;
   assign mem[165823:165792] = 32'b00000101011011010010101111011000;
   assign mem[165855:165824] = 32'b11111111110100111000011010001000;
   assign mem[165887:165856] = 32'b00000000001010010101001110110010;
   assign mem[165919:165888] = 32'b00000001000111011011101101011110;
   assign mem[165951:165920] = 32'b11111100110101010110101110101000;
   assign mem[165983:165952] = 32'b00000001001100000101100011111100;
   assign mem[166015:165984] = 32'b00000010011101100000010100001100;
   assign mem[166047:166016] = 32'b11111101110010101001110110011100;
   assign mem[166079:166048] = 32'b00000011110101010000000100010000;
   assign mem[166111:166080] = 32'b11111110101001110100000110101000;
   assign mem[166143:166112] = 32'b11111111111011110101110111011000;
   assign mem[166175:166144] = 32'b00000000001000101000001110001101;
   assign mem[166207:166176] = 32'b11111111110101100111100010110110;
   assign mem[166239:166208] = 32'b00000010100110000010110111010100;
   assign mem[166271:166240] = 32'b11111110010111100010100111011110;
   assign mem[166303:166272] = 32'b00000011011110110110010011011000;
   assign mem[166335:166304] = 32'b00000011000011111101001011111100;
   assign mem[166367:166336] = 32'b11111110001001000100011110100100;
   assign mem[166399:166368] = 32'b11111101101110100010011111110000;
   assign mem[166431:166400] = 32'b00000010101110001011111011011100;
   assign mem[166463:166432] = 32'b11111100110101001111011000110100;
   assign mem[166495:166464] = 32'b11111100100111100110100110101000;
   assign mem[166527:166496] = 32'b11111011000110110010110011110000;
   assign mem[166559:166528] = 32'b11110111001010101010001001000000;
   assign mem[166591:166560] = 32'b00000101011100101111001000111000;
   assign mem[166623:166592] = 32'b00000111001000011011110010001000;
   assign mem[166655:166624] = 32'b00000101101110111001011010001000;
   assign mem[166687:166656] = 32'b11110111111001111001100110100000;
   assign mem[166719:166688] = 32'b11111001100101100111010110011000;
   assign mem[166751:166720] = 32'b00000010011110011111001111010000;
   assign mem[166783:166752] = 32'b00000110111101111001111110011000;
   assign mem[166815:166784] = 32'b00001010100001000110001001000000;
   assign mem[166847:166816] = 32'b11110110010111000101011011010000;
   assign mem[166879:166848] = 32'b00000100001100111101001100100000;
   assign mem[166911:166880] = 32'b00000000001001011101010010001111;
   assign mem[166943:166912] = 32'b11111010100101001000000010100000;
   assign mem[166975:166944] = 32'b11110110111101011010101101000000;
   assign mem[167007:166976] = 32'b00000010000111011100001001111000;
   assign mem[167039:167008] = 32'b11111111101011110100110001101100;
   assign mem[167071:167040] = 32'b11111101110011001100100101101000;
   assign mem[167103:167072] = 32'b11111110101100101000111110011110;
   assign mem[167135:167104] = 32'b11111000011110010100110000110000;
   assign mem[167167:167136] = 32'b00000000110001110111100001010001;
   assign mem[167199:167168] = 32'b11110111000110011010001110000000;
   assign mem[167231:167200] = 32'b00000110001100000100000011000000;
   assign mem[167263:167232] = 32'b11111011111011001111111110111000;
   assign mem[167295:167264] = 32'b00000100000110110010101101101000;
   assign mem[167327:167296] = 32'b00000010101111111010111101111100;
   assign mem[167359:167328] = 32'b00000001001111110001010101000100;
   assign mem[167391:167360] = 32'b00000001010100001010011101011000;
   assign mem[167423:167392] = 32'b11111010000001001011100100110000;
   assign mem[167455:167424] = 32'b00000011101110011111001001100100;
   assign mem[167487:167456] = 32'b11111011000010111011110111110000;
   assign mem[167519:167488] = 32'b11111011111011110111110011001000;
   assign mem[167551:167520] = 32'b00000001001100110110111100111010;
   assign mem[167583:167552] = 32'b11111000111010110111111110101000;
   assign mem[167615:167584] = 32'b00000101111000101010000011101000;
   assign mem[167647:167616] = 32'b00000001001111110010100011100100;
   assign mem[167679:167648] = 32'b11111011111010010011010001000000;
   assign mem[167711:167680] = 32'b11111010000111000000111001011000;
   assign mem[167743:167712] = 32'b11110110001110000100111111100000;
   assign mem[167775:167744] = 32'b11110111101100111100001101000000;
   assign mem[167807:167776] = 32'b00001001111110100101111011100000;
   assign mem[167839:167808] = 32'b11111110000001011011001111111100;
   assign mem[167871:167840] = 32'b00000011010100111010101001000000;
   assign mem[167903:167872] = 32'b00000111101101000110111111000000;
   assign mem[167935:167904] = 32'b00000111111001011100100110001000;
   assign mem[167967:167936] = 32'b11111100100111000100110101011000;
   assign mem[167999:167968] = 32'b11101110010100001101110110100000;
   assign mem[168031:168000] = 32'b11111101001100001000111011010100;
   assign mem[168063:168032] = 32'b00000001100011011100100110000110;
   assign mem[168095:168064] = 32'b11111111001001010100000000011111;
   assign mem[168127:168096] = 32'b11111110111110111001110001100100;
   assign mem[168159:168128] = 32'b11111000001101111001110100111000;
   assign mem[168191:168160] = 32'b00000010000000010000010000011000;
   assign mem[168223:168192] = 32'b00000101110000110011001010001000;
   assign mem[168255:168224] = 32'b00000010111010000111100010100000;
   assign mem[168287:168256] = 32'b11111001110011011101001011011000;
   assign mem[168319:168288] = 32'b11111110110101011010000000010010;
   assign mem[168351:168320] = 32'b11111010101001110000100100010000;
   assign mem[168383:168352] = 32'b11111001011111111000101001111000;
   assign mem[168415:168384] = 32'b11110110111101100010101110110000;
   assign mem[168447:168416] = 32'b00001010000011110111001010110000;
   assign mem[168479:168448] = 32'b00000001010000011010001101011010;
   assign mem[168511:168480] = 32'b11111111010110011110110011010110;
   assign mem[168543:168512] = 32'b11111001000111001001111111001000;
   assign mem[168575:168544] = 32'b00000001110001011010000000111010;
   assign mem[168607:168576] = 32'b00000010001111101000110101011000;
   assign mem[168639:168608] = 32'b11111110100101111111100010111000;
   assign mem[168671:168640] = 32'b11111110001110111111101110100000;
   assign mem[168703:168672] = 32'b00000001110101001100000001001000;
   assign mem[168735:168704] = 32'b00000101000110001000001110111000;
   assign mem[168767:168736] = 32'b00000010101110100101100111111000;
   assign mem[168799:168768] = 32'b00000001001110011001010100101100;
   assign mem[168831:168800] = 32'b11101000010100100111101011000000;
   assign mem[168863:168832] = 32'b00000000111000011100011011100101;
   assign mem[168895:168864] = 32'b00000001100000110110100111100100;
   assign mem[168927:168896] = 32'b11111100111001010110011101010000;
   assign mem[168959:168928] = 32'b00000010101100001001001110000100;
   assign mem[168991:168960] = 32'b11111111101001101111111111111001;
   assign mem[169023:168992] = 32'b11111001010101101111100010110000;
   assign mem[169055:169024] = 32'b00000000111010010111111111011001;
   assign mem[169087:169056] = 32'b11111111011010100001000111001001;
   assign mem[169119:169088] = 32'b11111000010111111111111001111000;
   assign mem[169151:169120] = 32'b00001000100100010101100010010000;
   assign mem[169183:169152] = 32'b11111100110101010110111101011100;
   assign mem[169215:169184] = 32'b00000000011001010101010111010011;
   assign mem[169247:169216] = 32'b00000010000100011101001101110000;
   assign mem[169279:169248] = 32'b00000100100101001010101101101000;
   assign mem[169311:169280] = 32'b11111110101111110000100100101100;
   assign mem[169343:169312] = 32'b11111100101111001010000101100100;
   assign mem[169375:169344] = 32'b11111111010001111110111100010000;
   assign mem[169407:169376] = 32'b00000100000111000000010000111000;
   assign mem[169439:169408] = 32'b00000010000010110010001001110000;
   assign mem[169471:169440] = 32'b00000000101000010000110010001101;
   assign mem[169503:169472] = 32'b11110101001100101000110101010000;
   assign mem[169535:169504] = 32'b00001001110000111101111110000000;
   assign mem[169567:169536] = 32'b11111110010100101100000111100000;
   assign mem[169599:169568] = 32'b11111100101100011101001011011000;
   assign mem[169631:169600] = 32'b00000000111111010011100111101101;
   assign mem[169663:169632] = 32'b00000110010111110000111011111000;
   assign mem[169695:169664] = 32'b00000101010111011001010001100000;
   assign mem[169727:169696] = 32'b11111101110011110111010000111000;
   assign mem[169759:169728] = 32'b11110111001111111101101011010000;
   assign mem[169791:169760] = 32'b00001000000011111110001101010000;
   assign mem[169823:169792] = 32'b00001000001110111101101001100000;
   assign mem[169855:169824] = 32'b11111011101000001010110011010000;
   assign mem[169887:169856] = 32'b11110110100011111001011011000000;
   assign mem[169919:169888] = 32'b00000011000111001100000100001100;
   assign mem[169951:169920] = 32'b11101111000001001111101100000000;
   assign mem[169983:169952] = 32'b11101111000110100000100100100000;
   assign mem[170015:169984] = 32'b00000001111111101010101111010000;
   assign mem[170047:170016] = 32'b00000110101111001010111100000000;
   assign mem[170079:170048] = 32'b11110001000011100110111000110000;
   assign mem[170111:170080] = 32'b00000011001011001010101000011000;
   assign mem[170143:170112] = 32'b00000000100111100000000000111100;
   assign mem[170175:170144] = 32'b11111101110001011111000101001100;
   assign mem[170207:170176] = 32'b00001000111100011000110001100000;
   assign mem[170239:170208] = 32'b00000011110010110111011111000000;
   assign mem[170271:170240] = 32'b11111101000111001111110010111000;
   assign mem[170303:170272] = 32'b00001010001000001111011000110000;
   assign mem[170335:170304] = 32'b00000110011010001100100111110000;
   assign mem[170367:170336] = 32'b11111100101110101101110101010100;
   assign mem[170399:170368] = 32'b00000110100011011010100100000000;
   assign mem[170431:170400] = 32'b11110100101110111010000010110000;
   assign mem[170463:170432] = 32'b11110000011000101111000000010000;
   assign mem[170495:170464] = 32'b00000111000010101011100001010000;
   assign mem[170527:170496] = 32'b11111011110011001111100100000000;
   assign mem[170559:170528] = 32'b11111110101001010010100101000010;
   assign mem[170591:170560] = 32'b11111010101100010001110000100000;
   assign mem[170623:170592] = 32'b11111011000111101001101110111000;
   assign mem[170655:170624] = 32'b11111001110011111110100100010000;
   assign mem[170687:170656] = 32'b00000011011010011111000000000100;
   assign mem[170719:170688] = 32'b11110011101001011000100010000000;
   assign mem[170751:170720] = 32'b00000111100000111010010000000000;
   assign mem[170783:170752] = 32'b11111101101010010101101100101100;
   assign mem[170815:170784] = 32'b00000001010011010001100111101010;
   assign mem[170847:170816] = 32'b00000001011110001110111111100010;
   assign mem[170879:170848] = 32'b00000010110011110010010100111100;
   assign mem[170911:170880] = 32'b11111101000110000101100001011000;
   assign mem[170943:170912] = 32'b11111011000010000001011111101000;
   assign mem[170975:170944] = 32'b11111101100101000011010011101100;
   assign mem[171007:170976] = 32'b00001001111000111010111011010000;
   assign mem[171039:171008] = 32'b11111110101000101000111011100010;
   assign mem[171071:171040] = 32'b11111110000111010000000000010110;
   assign mem[171103:171072] = 32'b11111111110111011010010110101011;
   assign mem[171135:171104] = 32'b00000000010000000010110111011011;
   assign mem[171167:171136] = 32'b00000100101100000100010101110000;
   assign mem[171199:171168] = 32'b00000010011011000000110110001000;
   assign mem[171231:171200] = 32'b00001000101011011111000110100000;
   assign mem[171263:171232] = 32'b11111111001010110000101110001010;
   assign mem[171295:171264] = 32'b00000101011111111001110010010000;
   assign mem[171327:171296] = 32'b11111111010001111100110010110011;
   assign mem[171359:171328] = 32'b11111101101101111001100110111000;
   assign mem[171391:171360] = 32'b00000010001101101100001001011100;
   assign mem[171423:171392] = 32'b11101010101001001110001110100000;
   assign mem[171455:171424] = 32'b00000101000101011111001100000000;
   assign mem[171487:171456] = 32'b11111110111010101001111110001000;
   assign mem[171519:171488] = 32'b11111100010111101000010000000100;
   assign mem[171551:171520] = 32'b00000101010101011011110100000000;
   assign mem[171583:171552] = 32'b11111101011011100100001101111100;
   assign mem[171615:171584] = 32'b00000110111011011101001101001000;
   assign mem[171647:171616] = 32'b11111101111101100011100001110000;
   assign mem[171679:171648] = 32'b00000001101111011111110000101100;
   assign mem[171711:171680] = 32'b11110101000100111011111010110000;
   assign mem[171743:171712] = 32'b11101100000110011000110001100000;
   assign mem[171775:171744] = 32'b00000000011101000001000110010001;
   assign mem[171807:171776] = 32'b00000100001001111010000010000000;
   assign mem[171839:171808] = 32'b11111101011101111001111111001100;
   assign mem[171871:171840] = 32'b11111001011111100111110111011000;
   assign mem[171903:171872] = 32'b00000100000010000111111010100000;
   assign mem[171935:171904] = 32'b11111111101010101100111000010100;
   assign mem[171967:171936] = 32'b00000100110010001111001100111000;
   assign mem[171999:171968] = 32'b00000001111100101011010000010100;
   assign mem[172031:172000] = 32'b11110100101110101100100011000000;
   assign mem[172063:172032] = 32'b11111111011100110011011101101100;
   assign mem[172095:172064] = 32'b00000010110011000011011111010000;
   assign mem[172127:172096] = 32'b11111001111001000010101010110000;
   assign mem[172159:172128] = 32'b11111101100110011100101111011000;
   assign mem[172191:172160] = 32'b11111110111010111010111001110000;
   assign mem[172223:172192] = 32'b00000001001111011110100000000110;
   assign mem[172255:172224] = 32'b00000010100111010101000101000100;
   assign mem[172287:172256] = 32'b11111101010001110011010000110000;
   assign mem[172319:172288] = 32'b00000011100101111111101111111000;
   assign mem[172351:172320] = 32'b11110010000011101011001000100000;
   assign mem[172383:172352] = 32'b11111100010101110110101000010100;
   assign mem[172415:172384] = 32'b00000101110100010000100101111000;
   assign mem[172447:172416] = 32'b00000011100010110001010011100100;
   assign mem[172479:172448] = 32'b11111110001011111101000010111010;
   assign mem[172511:172480] = 32'b11110001100100010111100110100000;
   assign mem[172543:172512] = 32'b00010001111000100110011001100000;
   assign mem[172575:172544] = 32'b11111010101010000100101110110000;
   assign mem[172607:172576] = 32'b11110101011101110101100111100000;
   assign mem[172639:172608] = 32'b00000101011011100011101101111000;
   assign mem[172671:172640] = 32'b00001010001010101011111110010000;
   assign mem[172703:172672] = 32'b00001010010101000000011101110000;
   assign mem[172735:172704] = 32'b11111111101001010010111000100011;
   assign mem[172767:172736] = 32'b11111010010001100110111101101000;
   assign mem[172799:172768] = 32'b11110110001001000000010101000000;
   assign mem[172831:172800] = 32'b11111000111000111000110011111000;
   assign mem[172863:172832] = 32'b11101011000110100010011111000000;
   assign mem[172895:172864] = 32'b11111010001100110100110011001000;
   assign mem[172927:172896] = 32'b00000110010011100110110110010000;
   assign mem[172959:172928] = 32'b11110111011010110100101100100000;
   assign mem[172991:172960] = 32'b00000111110001110001011110011000;
   assign mem[173023:172992] = 32'b11111110110101101000100011011010;
   assign mem[173055:173024] = 32'b00000000101101100101100110011011;
   assign mem[173087:173056] = 32'b00001001010111110000101011100000;
   assign mem[173119:173088] = 32'b00000101110110110000001110111000;
   assign mem[173151:173120] = 32'b00000000101110000111000100111100;
   assign mem[173183:173152] = 32'b11111011011010100000110110100000;
   assign mem[173215:173184] = 32'b11111101100101001000011110001100;
   assign mem[173247:173216] = 32'b00000001001101001110011101010110;
   assign mem[173279:173248] = 32'b11110110111010001110010110000000;
   assign mem[173311:173280] = 32'b11111110101100100100011111010100;
   assign mem[173343:173312] = 32'b00000110001001101010110111101000;
   assign mem[173375:173344] = 32'b00000001010001011111101101010010;
   assign mem[173407:173376] = 32'b11111110111010001101000111110110;
   assign mem[173439:173408] = 32'b11111111111011101011101111001010;
   assign mem[173471:173440] = 32'b00000001010101011110110000110000;
   assign mem[173503:173472] = 32'b00000101100101100100011111011000;
   assign mem[173535:173504] = 32'b00000101100101101110011000101000;
   assign mem[173567:173536] = 32'b00000000001001010000011001110011;
   assign mem[173599:173568] = 32'b00000011100110010000011000101100;
   assign mem[173631:173600] = 32'b11110101101010100010001100110000;
   assign mem[173663:173632] = 32'b11111001001101010111001111101000;
   assign mem[173695:173664] = 32'b00000011011101100010000111101000;
   assign mem[173727:173696] = 32'b11111010111010100111101011000000;
   assign mem[173759:173728] = 32'b11111010111001111010001010000000;
   assign mem[173791:173760] = 32'b11111111111001000111101111010100;
   assign mem[173823:173792] = 32'b11110101010110010101100100000000;
   assign mem[173855:173824] = 32'b11111110110100011111011001110100;
   assign mem[173887:173856] = 32'b11111011111111101001100100001000;
   assign mem[173919:173888] = 32'b11101110001001001111111101100000;
   assign mem[173951:173920] = 32'b00001001000110100101110110000000;
   assign mem[173983:173952] = 32'b00000000011011000010101000001111;
   assign mem[174015:173984] = 32'b00000100000010111111000001101000;
   assign mem[174047:174016] = 32'b11111111100010110101101100101001;
   assign mem[174079:174048] = 32'b11111110000111011001001000111100;
   assign mem[174111:174080] = 32'b11111101001001010010010111100100;
   assign mem[174143:174112] = 32'b00000100000010100100100110001000;
   assign mem[174175:174144] = 32'b11110101110000100001011100010000;
   assign mem[174207:174176] = 32'b00000000000100111110011110001110;
   assign mem[174239:174208] = 32'b00000010011111001001011101001000;
   assign mem[174271:174240] = 32'b11111100101001011111110011100000;
   assign mem[174303:174272] = 32'b11111101100011100011110111011100;
   assign mem[174335:174304] = 32'b00000010100100001101000001110100;
   assign mem[174367:174336] = 32'b00000001000000111000100101011010;
   assign mem[174399:174368] = 32'b00000101000100101111100000011000;
   assign mem[174431:174400] = 32'b11111001000000010110010000000000;
   assign mem[174463:174432] = 32'b00000110111101110101001111001000;
   assign mem[174495:174464] = 32'b00000011101000110111101110010100;
   assign mem[174527:174496] = 32'b11110010111111100000111111000000;
   assign mem[174559:174528] = 32'b00000011100000111001011111111100;
   assign mem[174591:174560] = 32'b11111000111011011111000110110000;
   assign mem[174623:174592] = 32'b00000001101101011111111011011010;
   assign mem[174655:174624] = 32'b11111101011101000111100111011000;
   assign mem[174687:174656] = 32'b11111110010110110100100100000000;
   assign mem[174719:174688] = 32'b00000001010110110001000011101000;
   assign mem[174751:174720] = 32'b11111100101011010100110000111000;
   assign mem[174783:174752] = 32'b11110111001000011001011001100000;
   assign mem[174815:174784] = 32'b11111110001011000101111001100010;
   assign mem[174847:174816] = 32'b11111110001011010110011010110100;
   assign mem[174879:174848] = 32'b11110011000000101000111011110000;
   assign mem[174911:174880] = 32'b00000111101010000111001000100000;
   assign mem[174943:174912] = 32'b11111010001111110010101011111000;
   assign mem[174975:174944] = 32'b00000010011100111010111000010000;
   assign mem[175007:174976] = 32'b00000011011000100111001111010000;
   assign mem[175039:175008] = 32'b11111111111111101011001010101110;
   assign mem[175071:175040] = 32'b11110100101001000111111001010000;
   assign mem[175103:175072] = 32'b00000100110100111011001011111000;
   assign mem[175135:175104] = 32'b00000010000100001110000010111100;
   assign mem[175167:175136] = 32'b00000111001010001111100010011000;
   assign mem[175199:175168] = 32'b00000110110011100101011000111000;
   assign mem[175231:175200] = 32'b11111100011111011111111111011000;
   assign mem[175263:175232] = 32'b00000101010111101000100110100000;
   assign mem[175295:175264] = 32'b11111100110101000111000000001100;
   assign mem[175327:175296] = 32'b11111001111011010010101010100000;
   assign mem[175359:175328] = 32'b11110111000011010111010100010000;
   assign mem[175391:175360] = 32'b00000000010101111000100011011101;
   assign mem[175423:175392] = 32'b11111101111110101001111010101100;
   assign mem[175455:175424] = 32'b00000001010111001010011110010100;
   assign mem[175487:175456] = 32'b00000011110100011100101101010100;
   assign mem[175519:175488] = 32'b11110100110010100111011001010000;
   assign mem[175551:175520] = 32'b00000011000001111100011110011100;
   assign mem[175583:175552] = 32'b00000101011000111100010000001000;
   assign mem[175615:175584] = 32'b00000011100001110001100110100000;
   assign mem[175647:175616] = 32'b11111110001000011110001110101000;
   assign mem[175679:175648] = 32'b00000001111000011100101101010110;
   assign mem[175711:175680] = 32'b00000000011101001000110010100000;
   assign mem[175743:175712] = 32'b00000010010111000110110011010100;
   assign mem[175775:175744] = 32'b00000000111110001001101011010010;
   assign mem[175807:175776] = 32'b00000001001000010110001000000000;
   assign mem[175839:175808] = 32'b11111111000110111101110111100100;
   assign mem[175871:175840] = 32'b11111111111111101101001111010001;
   assign mem[175903:175872] = 32'b11111110111011100111011000001110;
   assign mem[175935:175904] = 32'b00000010111100000011001110011100;
   assign mem[175967:175936] = 32'b00000000010000000100101110011001;
   assign mem[175999:175968] = 32'b00000010110100111000001000110100;
   assign mem[176031:176000] = 32'b11111110010011001010110101101010;
   assign mem[176063:176032] = 32'b00001000111010111011100011100000;
   assign mem[176095:176064] = 32'b11111011110001110100111001100000;
   assign mem[176127:176096] = 32'b00000000101000000100101100000000;
   assign mem[176159:176128] = 32'b00000111111000101011011001001000;
   assign mem[176191:176160] = 32'b00000101101100111000000100100000;
   assign mem[176223:176192] = 32'b11110110100000000001010001010000;
   assign mem[176255:176224] = 32'b11111111101101000010100000110101;
   assign mem[176287:176256] = 32'b00000010100111001001000000101100;
   assign mem[176319:176288] = 32'b11111011110000000010001010001000;
   assign mem[176351:176320] = 32'b11110000011001001100100010110000;
   assign mem[176383:176352] = 32'b00001000000000001000100010010000;
   assign mem[176415:176384] = 32'b00000010000111110001101000010100;
   assign mem[176447:176416] = 32'b00000010100101100010000111111000;
   assign mem[176479:176448] = 32'b11110001100010000101100010100000;
   assign mem[176511:176480] = 32'b00000101100011101100011100000000;
   assign mem[176543:176512] = 32'b00000011011010000101000010001000;
   assign mem[176575:176544] = 32'b00000001001001011110001010110110;
   assign mem[176607:176576] = 32'b11111010101001000010110011000000;
   assign mem[176639:176608] = 32'b11111100101011111000010011001000;
   assign mem[176671:176640] = 32'b00000110110011001110011110001000;
   assign mem[176703:176672] = 32'b11111011101011101101110001111000;
   assign mem[176735:176704] = 32'b11111101101101011101000011100000;
   assign mem[176767:176736] = 32'b11111100110000000101000000111100;
   assign mem[176799:176768] = 32'b00000111101101010110110001100000;
   assign mem[176831:176800] = 32'b00000010000000010110111011111100;
   assign mem[176863:176832] = 32'b11111110110111111011101111111000;
   assign mem[176895:176864] = 32'b00000100100111101011001000101000;
   assign mem[176927:176896] = 32'b11111011000101010011101100000000;
   assign mem[176959:176928] = 32'b11111110001011011101110011100100;
   assign mem[176991:176960] = 32'b11111000101101110011000110111000;
   assign mem[177023:176992] = 32'b00000100111010011100011100011000;
   assign mem[177055:177024] = 32'b11111001001111000000001111001000;
   assign mem[177087:177056] = 32'b11111000001001111001000100001000;
   assign mem[177119:177088] = 32'b11111111101100100101100010010000;
   assign mem[177151:177120] = 32'b00001000111011000000000011010000;
   assign mem[177183:177152] = 32'b00000001100101100010011001011010;
   assign mem[177215:177184] = 32'b00000111011001111011110010000000;
   assign mem[177247:177216] = 32'b00000010111101110110010100101100;
   assign mem[177279:177248] = 32'b00000000100000111010111110000111;
   assign mem[177311:177280] = 32'b11111110011000001110001011011100;
   assign mem[177343:177312] = 32'b11110101001001010111001000000000;
   assign mem[177375:177344] = 32'b00000111010011110000001000100000;
   assign mem[177407:177376] = 32'b11110110011010101111100100100000;
   assign mem[177439:177408] = 32'b11110000010000110100111100000000;
   assign mem[177471:177440] = 32'b00000110101100010010101010100000;
   assign mem[177503:177472] = 32'b00001100000111010111110101000000;
   assign mem[177535:177504] = 32'b00000001100010000101100110101110;
   assign mem[177567:177536] = 32'b11110000111011011010100001010000;
   assign mem[177599:177568] = 32'b00000010010001000011001111101100;
   assign mem[177631:177600] = 32'b00000011001110011001101100101000;
   assign mem[177663:177632] = 32'b11111111011001011001001100110110;
   assign mem[177695:177664] = 32'b00000110101101011011000101110000;
   assign mem[177727:177696] = 32'b11111111111011110110010100100001;
   assign mem[177759:177728] = 32'b00000010000111000101010101010000;
   assign mem[177791:177760] = 32'b11101100011010101001101100100000;
   assign mem[177823:177792] = 32'b11110101111000100110110100110000;
   assign mem[177855:177824] = 32'b11111101110110010010000100101100;
   assign mem[177887:177856] = 32'b00000000010100001111011011100111;
   assign mem[177919:177888] = 32'b11111110101100000110001001100100;
   assign mem[177951:177920] = 32'b11111000010111001010110100100000;
   assign mem[177983:177952] = 32'b00001010101010110000111010100000;
   assign mem[178015:177984] = 32'b11111010100110010100011001100000;
   assign mem[178047:178016] = 32'b00001011110111110011011010000000;
   assign mem[178079:178048] = 32'b00000101001110001011001001001000;
   assign mem[178111:178080] = 32'b00000001011110111111101000001000;
   assign mem[178143:178112] = 32'b11101110111011101011100111100000;
   assign mem[178175:178144] = 32'b11101111100011001101011010000000;
   assign mem[178207:178176] = 32'b11111101111010000101111100100000;
   assign mem[178239:178208] = 32'b00000100100001000111010010010000;
   assign mem[178271:178240] = 32'b00000010001110011011000100011000;
   assign mem[178303:178272] = 32'b11111100100001110111100000101000;
   assign mem[178335:178304] = 32'b00000100111000110001011000001000;
   assign mem[178367:178336] = 32'b00000001010101101010001101110000;
   assign mem[178399:178368] = 32'b11111100000010111011010011111100;
   assign mem[178431:178400] = 32'b11110110000101100111001110110000;
   assign mem[178463:178432] = 32'b11111100011010000100110000000100;
   assign mem[178495:178464] = 32'b00000011011001111011111111000000;
   assign mem[178527:178496] = 32'b00000100101010001100011111101000;
   assign mem[178559:178528] = 32'b00000001111100000111000001010110;
   assign mem[178591:178560] = 32'b11111011101100101011111111000000;
   assign mem[178623:178592] = 32'b11111100100100001001010111111000;
   assign mem[178655:178624] = 32'b00000010000101101001001011101100;
   assign mem[178687:178656] = 32'b00000010001001010000000111111000;
   assign mem[178719:178688] = 32'b00000001000001001110100101101110;
   assign mem[178751:178720] = 32'b11111001011111110101000010100000;
   assign mem[178783:178752] = 32'b11111010111100010011010011111000;
   assign mem[178815:178784] = 32'b00000101010101101000010010011000;
   assign mem[178847:178816] = 32'b11111101101011101110101111000000;
   assign mem[178879:178848] = 32'b00000000010100010001110100010001;
   assign mem[178911:178880] = 32'b00000010010011010000101111011000;
   assign mem[178943:178912] = 32'b11111110111010010001111111010010;
   assign mem[178975:178944] = 32'b00000011101110010101111111100100;
   assign mem[179007:178976] = 32'b11111101000011100110101000101100;
   assign mem[179039:179008] = 32'b00000011001100001000100110110100;
   assign mem[179071:179040] = 32'b11111111101111101100011101011101;
   assign mem[179103:179072] = 32'b00000000101100110101001001110010;
   assign mem[179135:179104] = 32'b11111111011000111110101011000110;
   assign mem[179167:179136] = 32'b00000001111000001001010000010110;
   assign mem[179199:179168] = 32'b00000000000011010011001111100110;
   assign mem[179231:179200] = 32'b00000010000001111010100100001000;
   assign mem[179263:179232] = 32'b00000101111000110000110001010000;
   assign mem[179295:179264] = 32'b11110110011011000000101001000000;
   assign mem[179327:179296] = 32'b00000011100011100010110110110100;
   assign mem[179359:179328] = 32'b11110110011001011110010100000000;
   assign mem[179391:179360] = 32'b00000101000101000101001010101000;
   assign mem[179423:179392] = 32'b11111101001101101101100110111100;
   assign mem[179455:179424] = 32'b00000001010101011010011000100110;
   assign mem[179487:179456] = 32'b11111100001101010100011010001000;
   assign mem[179519:179488] = 32'b11111110111100010000100000001100;
   assign mem[179551:179520] = 32'b11110110111010100010001110110000;
   assign mem[179583:179552] = 32'b00001010010101111101000110000000;
   assign mem[179615:179584] = 32'b11111000001000011001111001101000;
   assign mem[179647:179616] = 32'b11110001111111001011011100100000;
   assign mem[179679:179648] = 32'b00001000001000010101100001000000;
   assign mem[179711:179680] = 32'b00000100111101100010011011110000;
   assign mem[179743:179712] = 32'b00001111010011010101100011000000;
   assign mem[179775:179744] = 32'b00000100010010010100101001100000;
   assign mem[179807:179776] = 32'b11111000100111010100011111110000;
   assign mem[179839:179808] = 32'b11111011010101101001010110101000;
   assign mem[179871:179840] = 32'b11111010111101001110011011011000;
   assign mem[179903:179872] = 32'b11110100110011010110101100100000;
   assign mem[179935:179904] = 32'b00000001011010011100100011111110;
   assign mem[179967:179936] = 32'b00000111101001100110101111001000;
   assign mem[179999:179968] = 32'b11111110111101111011001000010000;
   assign mem[180031:180000] = 32'b11110100110100001000101100110000;
   assign mem[180063:180032] = 32'b11111101100011011001110000110000;
   assign mem[180095:180064] = 32'b00000110110111001101111101011000;
   assign mem[180127:180096] = 32'b00000110000101101101100011011000;
   assign mem[180159:180128] = 32'b00000111001111111000001000010000;
   assign mem[180191:180160] = 32'b00000110110101100010101110111000;
   assign mem[180223:180192] = 32'b00001100011110100101110100100000;
   assign mem[180255:180224] = 32'b00001001001010111001010010010000;
   assign mem[180287:180256] = 32'b11110000010010011100011110000000;
   assign mem[180319:180288] = 32'b11111111001111010111100111100111;
   assign mem[180351:180320] = 32'b11101000100011000110011010000000;
   assign mem[180383:180352] = 32'b11111010111101110111110000010000;
   assign mem[180415:180384] = 32'b00000000110011111100000100110010;
   assign mem[180447:180416] = 32'b11111110010010000010010001100010;
   assign mem[180479:180448] = 32'b11111111011011000100000101001010;
   assign mem[180511:180480] = 32'b00000001000110100000110010010110;
   assign mem[180543:180512] = 32'b11110101010001000001110111000000;
   assign mem[180575:180544] = 32'b11111100111011001100001010100100;
   assign mem[180607:180576] = 32'b00000010001111110001000000100000;
   assign mem[180639:180608] = 32'b11111100100001111111010101111100;
   assign mem[180671:180640] = 32'b00001000101000100010000010100000;
   assign mem[180703:180672] = 32'b11110111111111100000010101100000;
   assign mem[180735:180704] = 32'b00000100000101110010010000001000;
   assign mem[180767:180736] = 32'b11111110010010000110111110010110;
   assign mem[180799:180768] = 32'b00000001101011101011010001011100;
   assign mem[180831:180800] = 32'b11111101011011000100011010100000;
   assign mem[180863:180832] = 32'b11110110110001111100110000000000;
   assign mem[180895:180864] = 32'b11111100100101001100010111111000;
   assign mem[180927:180896] = 32'b00001000100100001011000011010000;
   assign mem[180959:180928] = 32'b11110010010010111100101010110000;
   assign mem[180991:180960] = 32'b00001001000101011000000001110000;
   assign mem[181023:180992] = 32'b11111100111101001110000110011100;
   assign mem[181055:181024] = 32'b00000101010011011101010111001000;
   assign mem[181087:181056] = 32'b00000011001110101111001010001000;
   assign mem[181119:181088] = 32'b11111101010101111111000000011100;
   assign mem[181151:181120] = 32'b11111101000001111001000001100100;
   assign mem[181183:181152] = 32'b00000000001111100101001011001101;
   assign mem[181215:181184] = 32'b11111010100000011011111111101000;
   assign mem[181247:181216] = 32'b11111111110100000110001010010100;
   assign mem[181279:181248] = 32'b11111010010101111110101001100000;
   assign mem[181311:181280] = 32'b00000110110101100100100001100000;
   assign mem[181343:181312] = 32'b00000100111000100010101001011000;
   assign mem[181375:181344] = 32'b00000110111110100000110101110000;
   assign mem[181407:181376] = 32'b11111001011110101110001111011000;
   assign mem[181439:181408] = 32'b11111001000001111110101011100000;
   assign mem[181471:181440] = 32'b00000110111010101110101111100000;
   assign mem[181503:181472] = 32'b11111101110011110110100110010000;
   assign mem[181535:181504] = 32'b00000001100111010101100010010100;
   assign mem[181567:181536] = 32'b00000000010010011100011000100110;
   assign mem[181599:181568] = 32'b00000111101101010001001000101000;
   assign mem[181631:181600] = 32'b11110000110110011000011111110000;
   assign mem[181663:181632] = 32'b00000011111010011010000011001000;
   assign mem[181695:181664] = 32'b00000001000010000011101111011010;
   assign mem[181727:181696] = 32'b11111100011000010000010001100000;
   assign mem[181759:181728] = 32'b11111100101111000101011100110100;
   assign mem[181791:181760] = 32'b00000101000000100000001111111000;
   assign mem[181823:181792] = 32'b00000110011001001100110000001000;
   assign mem[181855:181824] = 32'b00000110011101101111100110010000;
   assign mem[181887:181856] = 32'b00000111001100000111101100100000;
   assign mem[181919:181888] = 32'b11111011101110001100011111000000;
   assign mem[181951:181920] = 32'b11101111010111110010100011100000;
   assign mem[181983:181952] = 32'b11110110100000100110111110110000;
   assign mem[182015:181984] = 32'b00000010101000101000011000001100;
   assign mem[182047:182016] = 32'b11111101011111100001111011011100;
   assign mem[182079:182048] = 32'b00000110111110010101000110100000;
   assign mem[182111:182080] = 32'b11111110111010101110110001100000;
   assign mem[182143:182112] = 32'b11110000001010110010000111100000;
   assign mem[182175:182144] = 32'b00000100010111101101001010011000;
   assign mem[182207:182176] = 32'b00000001011101011010001111100100;
   assign mem[182239:182208] = 32'b11111000110101010001111011110000;
   assign mem[182271:182240] = 32'b11111101111100001011000110010000;
   assign mem[182303:182272] = 32'b11111110010001101100011001001000;
   assign mem[182335:182304] = 32'b00000100100111110001010111110000;
   assign mem[182367:182336] = 32'b11111110101101110001000101010110;
   assign mem[182399:182368] = 32'b00000000001000001000101111111000;
   assign mem[182431:182400] = 32'b00000110101010000010011001011000;
   assign mem[182463:182432] = 32'b11111110100110000101111100100000;
   assign mem[182495:182464] = 32'b00001001100001000001110000000000;
   assign mem[182527:182496] = 32'b11111110001110001010011110110000;
   assign mem[182559:182528] = 32'b11111101110100101110100011100000;
   assign mem[182591:182560] = 32'b11111100000101111010001001101000;
   assign mem[182623:182592] = 32'b11111101110000000101011101010100;
   assign mem[182655:182624] = 32'b00000001000111101101000010101100;
   assign mem[182687:182656] = 32'b11111000011000101010001010010000;
   assign mem[182719:182688] = 32'b00000010010010101000100111111000;
   assign mem[182751:182720] = 32'b00000111011100111001100000000000;
   assign mem[182783:182752] = 32'b11111101010010010100010111011100;
   assign mem[182815:182784] = 32'b00000001010000100111011001111010;
   assign mem[182847:182816] = 32'b00000010101110100101010000100100;
   assign mem[182879:182848] = 32'b11111111010001010000000101100001;
   assign mem[182911:182880] = 32'b11111010011101000101000110111000;
   assign mem[182943:182912] = 32'b11110101000110100100100010100000;
   assign mem[182975:182944] = 32'b11111111101011010100111000010001;
   assign mem[183007:182976] = 32'b00000010110101111111111011010000;
   assign mem[183039:183008] = 32'b00000100011111010010110110100000;
   assign mem[183071:183040] = 32'b11111101101101000010110001000000;
   assign mem[183103:183072] = 32'b00010000011100010110000111000000;
   assign mem[183135:183104] = 32'b11110111001000110010010110010000;
   assign mem[183167:183136] = 32'b11110101101010111101101001010000;
   assign mem[183199:183168] = 32'b11111110100010110000111000100010;
   assign mem[183231:183200] = 32'b00000110011110100000111010000000;
   assign mem[183263:183232] = 32'b00001010000100001000001011100000;
   assign mem[183295:183264] = 32'b00000110000001100100001110000000;
   assign mem[183327:183296] = 32'b11111000010101100000111100011000;
   assign mem[183359:183328] = 32'b11111100110100010001101101110000;
   assign mem[183391:183360] = 32'b11111110100101011111100101011110;
   assign mem[183423:183392] = 32'b00010000011101001111011011000000;
   assign mem[183455:183424] = 32'b11110111101010100110100010000000;
   assign mem[183487:183456] = 32'b11110001010010110101111111100000;
   assign mem[183519:183488] = 32'b00000111101101110110011111011000;
   assign mem[183551:183520] = 32'b00000011110100100101001011110000;
   assign mem[183583:183552] = 32'b00001001110101101000011101100000;
   assign mem[183615:183584] = 32'b11111111100011101010110110101100;
   assign mem[183647:183616] = 32'b11111001100000011100011111010000;
   assign mem[183679:183648] = 32'b11111001111101010110010111101000;
   assign mem[183711:183680] = 32'b00000000010001001110011010111101;
   assign mem[183743:183712] = 32'b00001100111100011101100100010000;
   assign mem[183775:183744] = 32'b00000110001111110001110111010000;
   assign mem[183807:183776] = 32'b11100101001010001000110000100000;
   assign mem[183839:183808] = 32'b00001101000000010100010001110000;
   assign mem[183871:183840] = 32'b11101110000010111111101110100000;
   assign mem[183903:183872] = 32'b11111111001001110101110110000100;
   assign mem[183935:183904] = 32'b11110010110011001100101001000000;
   assign mem[183967:183936] = 32'b11110111010110010101100110000000;
   assign mem[183999:183968] = 32'b11110111110011010110100101000000;
   assign mem[184031:184000] = 32'b11111001101011110110010101100000;
   assign mem[184063:184032] = 32'b00001001101100001011110101110000;
   assign mem[184095:184064] = 32'b11111111001000011101110110010110;
   assign mem[184127:184096] = 32'b00000001011110100001010010111100;
   assign mem[184159:184128] = 32'b00001001110100100010110000000000;
   assign mem[184191:184160] = 32'b11101111001011011011100111100000;
   assign mem[184223:184192] = 32'b11111100000111000101100110111000;
   assign mem[184255:184224] = 32'b11111111000100100111000010000101;
   assign mem[184287:184256] = 32'b00000100100011010010000001111000;
   assign mem[184319:184288] = 32'b11111110111111010101011100000010;
   assign mem[184351:184320] = 32'b11111101010001000010100000110100;
   assign mem[184383:184352] = 32'b11111101001111010100111111111000;
   assign mem[184415:184384] = 32'b11111101001001101110111101100100;
   assign mem[184447:184416] = 32'b00000010011110010010110110001000;
   assign mem[184479:184448] = 32'b00001111011111000100011110110000;
   assign mem[184511:184480] = 32'b11111111100011100010111001001101;
   assign mem[184543:184512] = 32'b00001010101110000100001100110000;
   assign mem[184575:184544] = 32'b11110100010110000111110100010000;
   assign mem[184607:184576] = 32'b00000000110101000100100010110011;
   assign mem[184639:184608] = 32'b11101111100001111110001101000000;
   assign mem[184671:184640] = 32'b00000011010000001110111000000000;
   assign mem[184703:184672] = 32'b11111011000111110100001101010000;
   assign mem[184735:184704] = 32'b11111111011101000101011010000111;
   assign mem[184767:184736] = 32'b11111111100011010001010100000001;
   assign mem[184799:184768] = 32'b00000001010101110110001101100110;
   assign mem[184831:184800] = 32'b11110101010010010110000110110000;
   assign mem[184863:184832] = 32'b11111101100111001111010000101000;
   assign mem[184895:184864] = 32'b00000000100100100101010011110111;
   assign mem[184927:184896] = 32'b00000001010011111101100001000110;
   assign mem[184959:184928] = 32'b11111111111100101100100011011011;
   assign mem[184991:184960] = 32'b00001000100010100010011100110000;
   assign mem[185023:184992] = 32'b11111010010100010111010110010000;
   assign mem[185055:185024] = 32'b11111100100010110010110010101000;
   assign mem[185087:185056] = 32'b11111100110101100011110000000000;
   assign mem[185119:185088] = 32'b11110010011110010101111001100000;
   assign mem[185151:185120] = 32'b11111100001010111001000001010000;
   assign mem[185183:185152] = 32'b00000001100001101100110001100110;
   assign mem[185215:185184] = 32'b11111110001000111111110100011010;
   assign mem[185247:185216] = 32'b00001001011011001011100011000000;
   assign mem[185279:185248] = 32'b00000100100001001000111110000000;
   assign mem[185311:185280] = 32'b00000100000010010010100000101000;
   assign mem[185343:185312] = 32'b11110010000000100000110001000000;
   assign mem[185375:185344] = 32'b11110101101111110111111000000000;
   assign mem[185407:185376] = 32'b11110010011100001100101011100000;
   assign mem[185439:185408] = 32'b11110000000101010011100101010000;
   assign mem[185471:185440] = 32'b00001110001010011110110110000000;
   assign mem[185503:185472] = 32'b00000010100101101000110011110100;
   assign mem[185535:185504] = 32'b11101101101101111111110011100000;
   assign mem[185567:185536] = 32'b00000100011110010001101000001000;
   assign mem[185599:185568] = 32'b00000110011100101110100010000000;
   assign mem[185631:185600] = 32'b11110010000100101000111010010000;
   assign mem[185663:185632] = 32'b11111010101011101100110100111000;
   assign mem[185695:185664] = 32'b11101001000100001110100001000000;
   assign mem[185727:185696] = 32'b11110001001111010110010101110000;
   assign mem[185759:185728] = 32'b11111100000110110110101110100000;
   assign mem[185791:185760] = 32'b00001100000111010101110010100000;
   assign mem[185823:185792] = 32'b00010001000001011011110111000000;
   assign mem[185855:185824] = 32'b11111101100010001111000101000000;
   assign mem[185887:185856] = 32'b00000000000100110000110111011010;
   assign mem[185919:185888] = 32'b11110111000000110001101100000000;
   assign mem[185951:185920] = 32'b11111101101101000011110111111100;
   assign mem[185983:185952] = 32'b00000110001100101001011100000000;
   assign mem[186015:185984] = 32'b00000000011001101110000010100101;
   assign mem[186047:186016] = 32'b00000111001100000101110001110000;
   assign mem[186079:186048] = 32'b00001001000000111011101001000000;
   assign mem[186111:186080] = 32'b11110010001011001110100001100000;
   assign mem[186143:186112] = 32'b00000001000001001010010110110010;
   assign mem[186175:186144] = 32'b11111000110101000001101011001000;
   assign mem[186207:186176] = 32'b00000010000100011011000010100100;
   assign mem[186239:186208] = 32'b11111011100100100000110001110000;
   assign mem[186271:186240] = 32'b11110101101101000110110101000000;
   assign mem[186303:186272] = 32'b11111111110001010110000011000110;
   assign mem[186335:186304] = 32'b11111011100111010000001001111000;
   assign mem[186367:186336] = 32'b00000100001000111011101010110000;
   assign mem[186399:186368] = 32'b00000000001000011000101100110101;
   assign mem[186431:186400] = 32'b11111101000110110101000101100000;
   assign mem[186463:186432] = 32'b11111111101010011111111000001110;
   assign mem[186495:186464] = 32'b11111111100010101100000110111111;
   assign mem[186527:186496] = 32'b00000000101000001000010110101111;
   assign mem[186559:186528] = 32'b00000000110000101101100110101010;
   assign mem[186591:186560] = 32'b11110010001111001000010101010000;
   assign mem[186623:186592] = 32'b11111111110100101010100101011011;
   assign mem[186655:186624] = 32'b11111111010011100010100101010001;
   assign mem[186687:186656] = 32'b00000010101100100101011011100000;
   assign mem[186719:186688] = 32'b00000110001011011101101101010000;
   assign mem[186751:186720] = 32'b00000010001000111001010000010100;
   assign mem[186783:186752] = 32'b11111101101100000010000111011100;
   assign mem[186815:186784] = 32'b00000111101100000111111010000000;
   assign mem[186847:186816] = 32'b00000000110101000001000100000111;
   assign mem[186879:186848] = 32'b11110111101000011000000000100000;
   assign mem[186911:186880] = 32'b00000000010110001010001101001001;
   assign mem[186943:186912] = 32'b11111010110101101010101010100000;
   assign mem[186975:186944] = 32'b11111110000000110100001110000110;
   assign mem[187007:186976] = 32'b11111100101110100011010011101000;
   assign mem[187039:187008] = 32'b11111100101110011111100111110100;
   assign mem[187071:187040] = 32'b00000000000111110100101101011111;
   assign mem[187103:187072] = 32'b00001011000100110001100010100000;
   assign mem[187135:187104] = 32'b00000011111111010001100111011000;
   assign mem[187167:187136] = 32'b11111011001011011001010100111000;
   assign mem[187199:187168] = 32'b11111010101100101111000111101000;
   assign mem[187231:187200] = 32'b11111110111010100001000001110000;
   assign mem[187263:187232] = 32'b00001001010011100100001001100000;
   assign mem[187295:187264] = 32'b11111110111110011111001111010010;
   assign mem[187327:187296] = 32'b00000000001111011110111000100100;
   assign mem[187359:187328] = 32'b00000001011000100011000101110000;
   assign mem[187391:187360] = 32'b00000000011101000101001101001010;
   assign mem[187423:187392] = 32'b11111011001001110111110001011000;
   assign mem[187455:187424] = 32'b00000011000111010110000001110000;
   assign mem[187487:187456] = 32'b11111000000010010010110100010000;
   assign mem[187519:187488] = 32'b11101100100011011001000101000000;
   assign mem[187551:187520] = 32'b11111000110011001101110100010000;
   assign mem[187583:187552] = 32'b11110010101100100100000111010000;
   assign mem[187615:187584] = 32'b11101101010110111111000111100000;
   assign mem[187647:187616] = 32'b11110011001111000001001010010000;
   assign mem[187679:187648] = 32'b00000001010100100110101011000010;
   assign mem[187711:187680] = 32'b00001010101111011010100011010000;
   assign mem[187743:187712] = 32'b11111011101101000110001111110000;
   assign mem[187775:187744] = 32'b00000000101011000101101010100001;
   assign mem[187807:187776] = 32'b00000100001010110011101101101000;
   assign mem[187839:187808] = 32'b11111101100111000000010111011000;
   assign mem[187871:187840] = 32'b00001001111001100110011110110000;
   assign mem[187903:187872] = 32'b11110111101110110100000011100000;
   assign mem[187935:187904] = 32'b11111101000001111110001010110100;
   assign mem[187967:187936] = 32'b11110000110100011001111101010000;
   assign mem[187999:187968] = 32'b11111001011000100001001101100000;
   assign mem[188031:188000] = 32'b11111111011111111010110001001001;
   assign mem[188063:188032] = 32'b00000011111011110001010111111000;
   assign mem[188095:188064] = 32'b11111101111101000111010001110000;
   assign mem[188127:188096] = 32'b00000111010101111010100110101000;
   assign mem[188159:188128] = 32'b00000011111011000010010010111000;
   assign mem[188191:188160] = 32'b11111010001110011110101001110000;
   assign mem[188223:188192] = 32'b11110110111101011001001111100000;
   assign mem[188255:188224] = 32'b00000001010001000110000100000100;
   assign mem[188287:188256] = 32'b00000111011011001111011010111000;
   assign mem[188319:188288] = 32'b00000111100000011000000110110000;
   assign mem[188351:188320] = 32'b00000110001000010000011110010000;
   assign mem[188383:188352] = 32'b00000101100110111101001010011000;
   assign mem[188415:188384] = 32'b00000000111011011101011001011010;
   assign mem[188447:188416] = 32'b11111101010000010100010011011000;
   assign mem[188479:188448] = 32'b11101101000110000111000110000000;
   assign mem[188511:188480] = 32'b00000010100001101010110101101000;
   assign mem[188543:188512] = 32'b11110101100010001111010000100000;
   assign mem[188575:188544] = 32'b11111100000001011000011111000000;
   assign mem[188607:188576] = 32'b11111110001110001010100001011100;
   assign mem[188639:188608] = 32'b11111001010111011001011011100000;
   assign mem[188671:188640] = 32'b11111011111000011100001000100000;
   assign mem[188703:188672] = 32'b00001010100011010001000000000000;
   assign mem[188735:188704] = 32'b00000000001011010011101010000010;
   assign mem[188767:188736] = 32'b00000010111001110011010110110000;
   assign mem[188799:188768] = 32'b11111111001010101000100111011100;
   assign mem[188831:188800] = 32'b00000000000001100001101100110111;
   assign mem[188863:188832] = 32'b00000110000101010011011111001000;
   assign mem[188895:188864] = 32'b11111011101010101011100000100000;
   assign mem[188927:188896] = 32'b00001000110011010001110101100000;
   assign mem[188959:188928] = 32'b00000101101111011011111011001000;
   assign mem[188991:188960] = 32'b00000111111111010111011001000000;
   assign mem[189023:188992] = 32'b11111101100110101101011011010000;
   assign mem[189055:189024] = 32'b11111101111111000100011110011100;
   assign mem[189087:189056] = 32'b11111011000010110001101000001000;
   assign mem[189119:189088] = 32'b11111011110111111100110110100000;
   assign mem[189151:189120] = 32'b00000101011110011000010000100000;
   assign mem[189183:189152] = 32'b11111100010111111010101100001100;
   assign mem[189215:189184] = 32'b00001001100000001011001110010000;
   assign mem[189247:189216] = 32'b11111100110000100010100100111100;
   assign mem[189279:189248] = 32'b00001000110001110111010011110000;
   assign mem[189311:189280] = 32'b11101010011001111001011100100000;
   assign mem[189343:189312] = 32'b11110100010010011011001001110000;
   assign mem[189375:189344] = 32'b11111000000010011100010001010000;
   assign mem[189407:189376] = 32'b00001000100001111110100010100000;
   assign mem[189439:189408] = 32'b11110100110100010110001101010000;
   assign mem[189471:189440] = 32'b11110110000110011111110011000000;
   assign mem[189503:189472] = 32'b11111100000010100011111010001100;
   assign mem[189535:189504] = 32'b11110011111100110010001001110000;
   assign mem[189567:189536] = 32'b11111010010010100100111111011000;
   assign mem[189599:189568] = 32'b00000010101010011100100000001100;
   assign mem[189631:189600] = 32'b00001110000011101110010101010000;
   assign mem[189663:189632] = 32'b00000000101110101110111110100001;
   assign mem[189695:189664] = 32'b00001100001111101111001101100000;
   assign mem[189727:189696] = 32'b11111111110010000100011010100111;
   assign mem[189759:189728] = 32'b11111100010100001111101100111000;
   assign mem[189791:189760] = 32'b00000100100001011100111011001000;
   assign mem[189823:189792] = 32'b11111100001010000010100011011100;
   assign mem[189855:189824] = 32'b11111010111000011101011100011000;
   assign mem[189887:189856] = 32'b11111011000011101001011010000000;
   assign mem[189919:189888] = 32'b11110101000111100010100001000000;
   assign mem[189951:189920] = 32'b00000100111100010010110000100000;
   assign mem[189983:189952] = 32'b11111110100011001010000110011000;
   assign mem[190015:189984] = 32'b00000101110000100111101100000000;
   assign mem[190047:190016] = 32'b00000100110111010110001110111000;
   assign mem[190079:190048] = 32'b11111110110111010011010111111110;
   assign mem[190111:190080] = 32'b11111011111000111011010111010000;
   assign mem[190143:190112] = 32'b11110100110010010010110010100000;
   assign mem[190175:190144] = 32'b11111010111101111111011000101000;
   assign mem[190207:190176] = 32'b11111100101101001111101000111000;
   assign mem[190239:190208] = 32'b11111111100010110000110101100100;
   assign mem[190271:190240] = 32'b00001000100011010110010000000000;
   assign mem[190303:190272] = 32'b00000111001111111000111110110000;
   assign mem[190335:190304] = 32'b11111001011000011010111111101000;
   assign mem[190367:190336] = 32'b11111110101001100101011101001010;
   assign mem[190399:190368] = 32'b00000101010011010111110111010000;
   assign mem[190431:190400] = 32'b11111001111001010001001101001000;
   assign mem[190463:190432] = 32'b11101010010111010000000101100000;
   assign mem[190495:190464] = 32'b11111100010001011110000110011100;
   assign mem[190527:190496] = 32'b00000101101011011101001011001000;
   assign mem[190559:190528] = 32'b11111000011101101101100100100000;
   assign mem[190591:190560] = 32'b00000001000011000110111000000000;
   assign mem[190623:190592] = 32'b00001000111100010011000111110000;
   assign mem[190655:190624] = 32'b11111111110011111111001001111001;
   assign mem[190687:190656] = 32'b00000011001001100000100011000100;
   assign mem[190719:190688] = 32'b11111111100101010111001100000101;
   assign mem[190751:190720] = 32'b00000100001100110011011010111000;
   assign mem[190783:190752] = 32'b11111101011110011101111100001100;
   assign mem[190815:190784] = 32'b00000010010110111111100001000100;
   assign mem[190847:190816] = 32'b11111011000110111011010100100000;
   assign mem[190879:190848] = 32'b00001000101101000111010101100000;
   assign mem[190911:190880] = 32'b11110100100110010011101110100000;
   assign mem[190943:190912] = 32'b11110110110101001001011010010000;
   assign mem[190975:190944] = 32'b11110100111111100111100001110000;
   assign mem[191007:190976] = 32'b00000100110000101111100100010000;
   assign mem[191039:191008] = 32'b11111100000111001011110100010000;
   assign mem[191071:191040] = 32'b00000000011100011010000011011100;
   assign mem[191103:191072] = 32'b11110111101001001100001000100000;
   assign mem[191135:191104] = 32'b11111110101101100001110101001010;
   assign mem[191167:191136] = 32'b00000001101000011011100101011000;
   assign mem[191199:191168] = 32'b00000110001000010100111101001000;
   assign mem[191231:191200] = 32'b00000001000111101100100111100100;
   assign mem[191263:191232] = 32'b11111101101101110101110011111100;
   assign mem[191295:191264] = 32'b11111101010100101111101000001000;
   assign mem[191327:191296] = 32'b00000010111111111011001000100000;
   assign mem[191359:191328] = 32'b11111101110100010011101011111000;
   assign mem[191391:191360] = 32'b11110101111000010101100101010000;
   assign mem[191423:191392] = 32'b00000001101110010001011111100110;
   assign mem[191455:191424] = 32'b00000011011101100110010011001000;
   assign mem[191487:191456] = 32'b00000100110110111110010000100000;
   assign mem[191519:191488] = 32'b00000011000101100000111100111100;
   assign mem[191551:191520] = 32'b11101101100101010000010101000000;
   assign mem[191583:191552] = 32'b11110100101000101100101101100000;
   assign mem[191615:191584] = 32'b00000101100110100110100001101000;
   assign mem[191647:191616] = 32'b00000101100100111110110110000000;
   assign mem[191679:191648] = 32'b11111111110110000000101001101111;
   assign mem[191711:191680] = 32'b00000111001101001100100010010000;
   assign mem[191743:191712] = 32'b11111101111100001001111111100000;
   assign mem[191775:191744] = 32'b11111111100010110110101110100000;
   assign mem[191807:191776] = 32'b11111101001001000011010101000000;
   assign mem[191839:191808] = 32'b00000001110010110110111110011000;
   assign mem[191871:191840] = 32'b11110001000011110101110111010000;
   assign mem[191903:191872] = 32'b11110101101110110011011111110000;
   assign mem[191935:191904] = 32'b11111011110001111010101011000000;
   assign mem[191967:191936] = 32'b00000011100100100111000101000000;
   assign mem[191999:191968] = 32'b00000100000001101000010101000000;
   assign mem[192031:192000] = 32'b00001011001101101011001000110000;
   assign mem[192063:192032] = 32'b11111110110100110011101001101010;
   assign mem[192095:192064] = 32'b00000000011001100000001101010110;
   assign mem[192127:192096] = 32'b11110110110001110000100001010000;
   assign mem[192159:192128] = 32'b00000110110110011100101001111000;
   assign mem[192191:192160] = 32'b11101100000011000010101011100000;
   assign mem[192223:192192] = 32'b11111101001100101111101111010100;
   assign mem[192255:192224] = 32'b11111101000010101011110111100000;
   assign mem[192287:192256] = 32'b00000111011110111111011111001000;
   assign mem[192319:192288] = 32'b11111100110100100100101100010000;
   assign mem[192351:192320] = 32'b11111101010101111100011100110000;
   assign mem[192383:192352] = 32'b11111101110111001010111001010100;
   assign mem[192415:192384] = 32'b11111111000011100011010101110101;
   assign mem[192447:192416] = 32'b00000010001001100111010001000100;
   assign mem[192479:192448] = 32'b11111111100001101110011001000000;
   assign mem[192511:192480] = 32'b11111010011001111010000111001000;
   assign mem[192543:192512] = 32'b11111010110011101111110100011000;
   assign mem[192575:192544] = 32'b00000011001000101111110011100100;
   assign mem[192607:192576] = 32'b00000000011100011010010100001101;
   assign mem[192639:192608] = 32'b00000001100010001111111100100100;
   assign mem[192671:192640] = 32'b00000100000011000001101100010000;
   assign mem[192703:192672] = 32'b00000001001011101101110001101000;
   assign mem[192735:192704] = 32'b00000001001010011100111111001100;
   assign mem[192767:192736] = 32'b00000000110111001000100001101000;
   assign mem[192799:192768] = 32'b00000011000110110010000001110000;
   assign mem[192831:192800] = 32'b11110010111111000101010001110000;
   assign mem[192863:192832] = 32'b11101011000111010111010011100000;
   assign mem[192895:192864] = 32'b11111101010101111000110011010100;
   assign mem[192927:192896] = 32'b00000000100100010001100110111100;
   assign mem[192959:192928] = 32'b00000011011000101101101110101000;
   assign mem[192991:192960] = 32'b11100110011111100000011101000000;
   assign mem[193023:192992] = 32'b00001000101001000110100101110000;
   assign mem[193055:193024] = 32'b11110101111010111111110000100000;
   assign mem[193087:193056] = 32'b11111001111000011010000000001000;
   assign mem[193119:193088] = 32'b00000100000011011000001111001000;
   assign mem[193151:193120] = 32'b00001010000111100100011011110000;
   assign mem[193183:193152] = 32'b00000101001110101011001100100000;
   assign mem[193215:193184] = 32'b00001010110001100101011100000000;
   assign mem[193247:193216] = 32'b11111111000001001101101110111000;
   assign mem[193279:193248] = 32'b11101011100011000110000111100000;
   assign mem[193311:193280] = 32'b11110111111001100111110011100000;
   assign mem[193343:193312] = 32'b11111001011111011110001000000000;
   assign mem[193375:193344] = 32'b11111101010010011001110101100000;
   assign mem[193407:193376] = 32'b00000100011111100110010010010000;
   assign mem[193439:193408] = 32'b11111111100101011011101011010100;
   assign mem[193471:193440] = 32'b00000111000000100111100100101000;
   assign mem[193503:193472] = 32'b11110111111010110010001100100000;
   assign mem[193535:193504] = 32'b11111111110100000001010101010110;
   assign mem[193567:193536] = 32'b00000011011110101011000101000000;
   assign mem[193599:193568] = 32'b11111100110101110011111100110100;
   assign mem[193631:193600] = 32'b00000100000110111111010110010000;
   assign mem[193663:193632] = 32'b11110010110101101010100100110000;
   assign mem[193695:193664] = 32'b11111101011001111110010011001000;
   assign mem[193727:193696] = 32'b11111100001100110111110110010100;
   assign mem[193759:193728] = 32'b11110011100100000011100001100000;
   assign mem[193791:193760] = 32'b00000010110001011001001000001100;
   assign mem[193823:193792] = 32'b00001001101011110011100010110000;
   assign mem[193855:193824] = 32'b00000000110101000101000101100110;
   assign mem[193887:193856] = 32'b00000010000000101011100010001000;
   assign mem[193919:193888] = 32'b11111010110001001101111101001000;
   assign mem[193951:193920] = 32'b00000111001011100011001000000000;
   assign mem[193983:193952] = 32'b11110111001101000101011110000000;
   assign mem[194015:193984] = 32'b00000101110010010000000011011000;
   assign mem[194047:194016] = 32'b11111100110001101010000011110100;
   assign mem[194079:194048] = 32'b00000000010101010011100101111111;
   assign mem[194111:194080] = 32'b11110001001110110001111010110000;
   assign mem[194143:194112] = 32'b11101110000001001110100001000000;
   assign mem[194175:194144] = 32'b00000100001110111000011000010000;
   assign mem[194207:194176] = 32'b00000100111111110100001001011000;
   assign mem[194239:194208] = 32'b00000010001110100101111101011000;
   assign mem[194271:194240] = 32'b00000010100010001010011101000000;
   assign mem[194303:194272] = 32'b11111000111001111100100100010000;
   assign mem[194335:194304] = 32'b11101001001101001110010110000000;
   assign mem[194367:194336] = 32'b11111000011101010100111011100000;
   assign mem[194399:194368] = 32'b00000000000010110110100101101001;
   assign mem[194431:194400] = 32'b00001011011000010000110010100000;
   assign mem[194463:194432] = 32'b00000011101101010000010010011100;
   assign mem[194495:194464] = 32'b11111010011100111001001000111000;
   assign mem[194527:194496] = 32'b11111111110101100101010000000000;
   assign mem[194559:194528] = 32'b11111100111100101010100000111100;
   assign mem[194591:194560] = 32'b11111110011000101101110010010110;
   assign mem[194623:194592] = 32'b00000111111110101001110001011000;
   assign mem[194655:194624] = 32'b11110001010001010010000100100000;
   assign mem[194687:194656] = 32'b00000110000100111100000000110000;
   assign mem[194719:194688] = 32'b00000111111001000111110010100000;
   assign mem[194751:194720] = 32'b11111100111001000001110110111000;
   assign mem[194783:194752] = 32'b00000000000100100000001111101101;
   assign mem[194815:194784] = 32'b00001111001110101000110000110000;
   assign mem[194847:194816] = 32'b11111010100010101000110111001000;
   assign mem[194879:194848] = 32'b11111001100100100010100111110000;
   assign mem[194911:194880] = 32'b00000011110000011001000110010000;
   assign mem[194943:194912] = 32'b00001001010110100010000100100000;
   assign mem[194975:194944] = 32'b00000011101011010111001101110000;
   assign mem[195007:194976] = 32'b11110001111100101011000100110000;
   assign mem[195039:195008] = 32'b00000110011001111100011001110000;
   assign mem[195071:195040] = 32'b11111000100001111000111010010000;
   assign mem[195103:195072] = 32'b11111001011011010111101111010000;
   assign mem[195135:195104] = 32'b11110111110111111000111001010000;
   assign mem[195167:195136] = 32'b00000010101010100010111111011000;
   assign mem[195199:195168] = 32'b11110110010100001111001000010000;
   assign mem[195231:195200] = 32'b00000010111011000100110101100100;
   assign mem[195263:195232] = 32'b11111111011111010101101010011101;
   assign mem[195295:195264] = 32'b11111000001010110010110100011000;
   assign mem[195327:195296] = 32'b11111101000111000001110100010000;
   assign mem[195359:195328] = 32'b11111110001111000111011100110010;
   assign mem[195391:195360] = 32'b00001000101101100111000010000000;
   assign mem[195423:195392] = 32'b11111110010000111011001100011000;
   assign mem[195455:195424] = 32'b11110111100011100000100000010000;
   assign mem[195487:195456] = 32'b00000110001100010001001010011000;
   assign mem[195519:195488] = 32'b00000000100001110010100100010010;
   assign mem[195551:195520] = 32'b11110011110111011100100111000000;
   assign mem[195583:195552] = 32'b00000001110110001110101110110000;
   assign mem[195615:195584] = 32'b11111110010010011100010100010010;
   assign mem[195647:195616] = 32'b00000001111110100111111110010110;
   assign mem[195679:195648] = 32'b00000000100001001111000111011011;
   assign mem[195711:195680] = 32'b11111110011011000110010101100010;
   assign mem[195743:195712] = 32'b11111100010011111001010110110000;
   assign mem[195775:195744] = 32'b00000101101100011000101101100000;
   assign mem[195807:195776] = 32'b00000001100101100111111010011000;
   assign mem[195839:195808] = 32'b11111110110011100101110101011010;
   assign mem[195871:195840] = 32'b00000010010001010010010111111100;
   assign mem[195903:195872] = 32'b11110000000100010001110010110000;
   assign mem[195935:195904] = 32'b00000000100000101000110111001110;
   assign mem[195967:195936] = 32'b11111011000110000100100101010000;
   assign mem[195999:195968] = 32'b11111100101110100010011101111000;
   assign mem[196031:196000] = 32'b00000010111000010110101001011100;
   assign mem[196063:196032] = 32'b00001010000001101100000011100000;
   assign mem[196095:196064] = 32'b11111111010000100101011011110011;
   assign mem[196127:196096] = 32'b11111110001000111001000100011110;
   assign mem[196159:196128] = 32'b00000010011100111010000000000000;
   assign mem[196191:196160] = 32'b00000011000110101000000011100000;
   assign mem[196223:196192] = 32'b11111001011011100100010011001000;
   assign mem[196255:196224] = 32'b11111101101001001111100100110000;
   assign mem[196287:196256] = 32'b11111100000101100010111011111000;
   assign mem[196319:196288] = 32'b11111001111000111001001100101000;
   assign mem[196351:196320] = 32'b00000000111001111110111001011001;
   assign mem[196383:196352] = 32'b00000011110100001110000101000000;
   assign mem[196415:196384] = 32'b11111111010000011000000101011010;
   assign mem[196447:196416] = 32'b00000011111001101100010100000100;
   assign mem[196479:196448] = 32'b00000000100101010010110100110110;
   assign mem[196511:196480] = 32'b11111111001110101000001000010111;
   assign mem[196543:196512] = 32'b11111000000111110001110111101000;
   assign mem[196575:196544] = 32'b11111110110010000101100101010000;
   assign mem[196607:196576] = 32'b11111101101101000100000000101000;
   assign mem[196639:196608] = 32'b00000101010110101000010110001000;
   assign mem[196671:196640] = 32'b00001001000110011001000111110000;
   assign mem[196703:196672] = 32'b11111110101000000100010100100100;
   assign mem[196735:196704] = 32'b11111000110010101010100000001000;
   assign mem[196767:196736] = 32'b11111100100110111101101001010000;
   assign mem[196799:196768] = 32'b00000011110110101110110110011000;
   assign mem[196831:196800] = 32'b00000000100110011000000011001111;
   assign mem[196863:196832] = 32'b11110100010111110010101110110000;
   assign mem[196895:196864] = 32'b11111100010000001001110001011000;
   assign mem[196927:196896] = 32'b11100111001101001101001000100000;
   assign mem[196959:196928] = 32'b11110101011000101010111100100000;
   assign mem[196991:196960] = 32'b00001100001101010110010101100000;
   assign mem[197023:196992] = 32'b00001100101111001011101001100000;
   assign mem[197055:197024] = 32'b11110110111110010000011001110000;
   assign mem[197087:197056] = 32'b00000001101000001111001010010000;
   assign mem[197119:197088] = 32'b11111000011111101100101100011000;
   assign mem[197151:197120] = 32'b00001101110000010010000111010000;
   assign mem[197183:197152] = 32'b11110101011000001110111101100000;
   assign mem[197215:197184] = 32'b00000001111110011001001001000000;
   assign mem[197247:197216] = 32'b11111100001110100010010101110100;
   assign mem[197279:197248] = 32'b00000010010001010010001000001100;
   assign mem[197311:197280] = 32'b11111010101010001111010011111000;
   assign mem[197343:197312] = 32'b00000100001100100010000101111000;
   assign mem[197375:197344] = 32'b00000001001110101000011010101100;
   assign mem[197407:197376] = 32'b00000010001000101000100101000000;
   assign mem[197439:197408] = 32'b11111111001110111110101101111100;
   assign mem[197471:197440] = 32'b11110100010001110100011010100000;
   assign mem[197503:197472] = 32'b11111110100111111110110110001110;
   assign mem[197535:197504] = 32'b11101100100010110001011000100000;
   assign mem[197567:197536] = 32'b11111100011011011000011111111000;
   assign mem[197599:197568] = 32'b00000010001001100111111010111000;
   assign mem[197631:197600] = 32'b00001001001001111000101110110000;
   assign mem[197663:197632] = 32'b00000101000101111100101001010000;
   assign mem[197695:197664] = 32'b00000001101110010100100101000010;
   assign mem[197727:197696] = 32'b11111111101100000011000111111011;
   assign mem[197759:197728] = 32'b11111111111110111101101010001010;
   assign mem[197791:197760] = 32'b11111011100110110111100010110000;
   assign mem[197823:197792] = 32'b11110111111011000011110010000000;
   assign mem[197855:197824] = 32'b11110000001001100111100001100000;
   assign mem[197887:197856] = 32'b11101000000001001000000001100000;
   assign mem[197919:197888] = 32'b11110011100111100001100110100000;
   assign mem[197951:197920] = 32'b00001010111101110101000111110000;
   assign mem[197983:197952] = 32'b00010010111101110111111000000000;
   assign mem[198015:197984] = 32'b11110110110111100101001101100000;
   assign mem[198047:198016] = 32'b11110101000100011110001101000000;
   assign mem[198079:198048] = 32'b11111001001000111010100001111000;
   assign mem[198111:198080] = 32'b00000001110001000001000101101100;
   assign mem[198143:198112] = 32'b11111101000000100001101001111100;
   assign mem[198175:198144] = 32'b00000001001110101011011001111100;
   assign mem[198207:198176] = 32'b00000011000011011110011111001000;
   assign mem[198239:198208] = 32'b00000000101011000111001100101110;
   assign mem[198271:198240] = 32'b11110000011011111000011001010000;
   assign mem[198303:198272] = 32'b11111000111001000111001010100000;
   assign mem[198335:198304] = 32'b00000001001010010111000001010110;
   assign mem[198367:198336] = 32'b11111111100000100100100100110110;
   assign mem[198399:198368] = 32'b00000001111011001111111010110100;
   assign mem[198431:198400] = 32'b11111110101110000011101110010100;
   assign mem[198463:198432] = 32'b00000011110111000101111100111100;
   assign mem[198495:198464] = 32'b11110111101100110000100000010000;
   assign mem[198527:198496] = 32'b00000011001100001010111101010000;
   assign mem[198559:198528] = 32'b00000011010101000101111001000000;
   assign mem[198591:198560] = 32'b11111111000110110000011101000101;
   assign mem[198623:198592] = 32'b11111111000111000100011011001111;
   assign mem[198655:198624] = 32'b11111110011000011111000010110100;
   assign mem[198687:198656] = 32'b11111011110100111111111001000000;
   assign mem[198719:198688] = 32'b11111111010010100011111100110101;
   assign mem[198751:198720] = 32'b00000101100110001010010011111000;
   assign mem[198783:198752] = 32'b11111100010011100010100000001000;
   assign mem[198815:198784] = 32'b00000001000100101011110101010110;
   assign mem[198847:198816] = 32'b11111111100101010010010101101111;
   assign mem[198879:198848] = 32'b11110010101001101110110001110000;
   assign mem[198911:198880] = 32'b11110101001110000011101001100000;
   assign mem[198943:198912] = 32'b00000000100101100101011111100111;
   assign mem[198975:198944] = 32'b00000000111101000101101011010001;
   assign mem[199007:198976] = 32'b00000100011101000110001000011000;
   assign mem[199039:199008] = 32'b00000101110001101110001100000000;
   assign mem[199071:199040] = 32'b00001001101011010001000110110000;
   assign mem[199103:199072] = 32'b11101111001011100110111100000000;
   assign mem[199135:199104] = 32'b00000101001000111001101001000000;
   assign mem[199167:199136] = 32'b11110001101101100100101111000000;
   assign mem[199199:199168] = 32'b11110111111011101010100010010000;
   assign mem[199231:199200] = 32'b00000111011111110110110000010000;
   assign mem[199263:199232] = 32'b11111110100000100000101101000110;
   assign mem[199295:199264] = 32'b11110010110000001111000011000000;
   assign mem[199327:199296] = 32'b00000100101101001101110101011000;
   assign mem[199359:199328] = 32'b11111101101001010101001001101000;
   assign mem[199391:199360] = 32'b00000001110000001111011011111000;
   assign mem[199423:199392] = 32'b11111100011110111101110000011000;
   assign mem[199455:199424] = 32'b11111110100100100010011001111010;
   assign mem[199487:199456] = 32'b11111101000010101101000000000000;
   assign mem[199519:199488] = 32'b11111100100100011010011011001100;
   assign mem[199551:199520] = 32'b11111101010001101010000000000000;
   assign mem[199583:199552] = 32'b11111100110101101110010001001000;
   assign mem[199615:199584] = 32'b11111111011001110111110111010010;
   assign mem[199647:199616] = 32'b11111110100010100000111001010000;
   assign mem[199679:199648] = 32'b00000001001100101000000110010100;
   assign mem[199711:199680] = 32'b11111110010100000100111010010000;
   assign mem[199743:199712] = 32'b00000110100111101010000100111000;
   assign mem[199775:199744] = 32'b11110011111010000111001100110000;
   assign mem[199807:199776] = 32'b11111110011000101111110001000100;
   assign mem[199839:199808] = 32'b00000001000011011111010010001100;
   assign mem[199871:199840] = 32'b00001000101010011000001110110000;
   assign mem[199903:199872] = 32'b11111001110000110010010101100000;
   assign mem[199935:199904] = 32'b00000011110111101100011010001000;
   assign mem[199967:199936] = 32'b11111101000101110010000001001000;
   assign mem[199999:199968] = 32'b11111111100111001110011110000111;
   assign mem[200031:200000] = 32'b11111000111101110100000110010000;
   assign mem[200063:200032] = 32'b00000111001110001001010110110000;
   assign mem[200095:200064] = 32'b11111100001000010100000111110000;
   assign mem[200127:200096] = 32'b11110111010000100010011000010000;
   assign mem[200159:200128] = 32'b00001000001110001101001110110000;
   assign mem[200191:200160] = 32'b11111111011011100110100011101101;
   assign mem[200223:200192] = 32'b00000110100010001111100101100000;
   assign mem[200255:200224] = 32'b00000111001111000010001110001000;
   assign mem[200287:200256] = 32'b00000100010101000000001110100000;
   assign mem[200319:200288] = 32'b11101000111110001011101110100000;
   assign mem[200351:200320] = 32'b11111111000110110100110000110001;
   assign mem[200383:200352] = 32'b11111011111101100000010111011000;
   assign mem[200415:200384] = 32'b00000110000101000011100110101000;
   assign mem[200447:200416] = 32'b00001000101101000101000110010000;
   assign mem[200479:200448] = 32'b00000010000110111001100001010000;
   assign mem[200511:200480] = 32'b11101100101101100010111000000000;
   assign mem[200543:200512] = 32'b11111001010001101111110001100000;
   assign mem[200575:200544] = 32'b00000010011010110111011010000000;
   assign mem[200607:200576] = 32'b00000101001010010001100110111000;
   assign mem[200639:200608] = 32'b11111100111100111110101111001000;
   assign mem[200671:200640] = 32'b00000100010100101110101111010000;
   assign mem[200703:200672] = 32'b00000111001001001111001111010000;
   assign mem[200735:200704] = 32'b00000010010001101101100111001100;
   assign mem[200767:200736] = 32'b11111001111110010101001101001000;
   assign mem[200799:200768] = 32'b00000000110010101010001111011101;
   assign mem[200831:200800] = 32'b11101111010100010001111000000000;
   assign mem[200863:200832] = 32'b00000000101010100010100011010011;
   assign mem[200895:200864] = 32'b11111101110001111111010011110100;
   assign mem[200927:200896] = 32'b00000011111010100110100001111100;
   assign mem[200959:200928] = 32'b11110110001011000010000010010000;
   assign mem[200991:200960] = 32'b00000011100110101110110100010100;
   assign mem[201023:200992] = 32'b11111101101110111111001000011000;
   assign mem[201055:201024] = 32'b11110101011010100100011110010000;
   assign mem[201087:201056] = 32'b11110100000100110100001011100000;
   assign mem[201119:201088] = 32'b11111010000010111001111111011000;
   assign mem[201151:201120] = 32'b00001101011111011110100000110000;
   assign mem[201183:201152] = 32'b00000010101111101110110001101000;
   assign mem[201215:201184] = 32'b00000000011000001100000101110000;
   assign mem[201247:201216] = 32'b00000100010011100001101111011000;
   assign mem[201279:201248] = 32'b00000000111111000100011110011100;
   assign mem[201311:201280] = 32'b11111110010011011000000110101110;
   assign mem[201343:201312] = 32'b11110011001111101100011001110000;
   assign mem[201375:201344] = 32'b11110111001100000011110100010000;
   assign mem[201407:201376] = 32'b11111001101010001011100111101000;
   assign mem[201439:201408] = 32'b11110111011010011011110111000000;
   assign mem[201471:201440] = 32'b00001011100111011100011110110000;
   assign mem[201503:201472] = 32'b11111100110110111110000111100100;
   assign mem[201535:201504] = 32'b11111101011101100111101011000000;
   assign mem[201567:201536] = 32'b00000110110100100111010000010000;
   assign mem[201599:201568] = 32'b11111011001000011000101111110000;
   assign mem[201631:201600] = 32'b11110111111011010010001111010000;
   assign mem[201663:201632] = 32'b00000011000111110111110111101000;
   assign mem[201695:201664] = 32'b11101111011001011010001111000000;
   assign mem[201727:201696] = 32'b00000100000000110110101101000000;
   assign mem[201759:201728] = 32'b00000010001000000110010010100100;
   assign mem[201791:201760] = 32'b00001001100010100100010001100000;
   assign mem[201823:201792] = 32'b11111111111011011110010100010010;
   assign mem[201855:201824] = 32'b00000101100111110110011110001000;
   assign mem[201887:201856] = 32'b00000011101101010100000011101100;
   assign mem[201919:201888] = 32'b11111001010010010010111000110000;
   assign mem[201951:201920] = 32'b11111101000011101100001111110100;
   assign mem[201983:201952] = 32'b00000001100000111101011000111000;
   assign mem[202015:201984] = 32'b00000000101000100101010001001001;
   assign mem[202047:202016] = 32'b00000110000010000010000100001000;
   assign mem[202079:202048] = 32'b11111111011101001111101110100010;
   assign mem[202111:202080] = 32'b11110000101001111011110011010000;
   assign mem[202143:202112] = 32'b11111000101111010100110101100000;
   assign mem[202175:202144] = 32'b00000011001010000011111001011100;
   assign mem[202207:202176] = 32'b00000100101101100101000011000000;
   assign mem[202239:202208] = 32'b11111011000000100101010000100000;
   assign mem[202271:202240] = 32'b00000010011101111110110100101100;
   assign mem[202303:202272] = 32'b00000000001100011101111100101111;
   assign mem[202335:202304] = 32'b00000001011000001101111000110110;
   assign mem[202367:202336] = 32'b00000101101111010001110001010000;
   assign mem[202399:202368] = 32'b11111100111100000100110011001100;
   assign mem[202431:202400] = 32'b11110000101010100100100100010000;
   assign mem[202463:202432] = 32'b11110000110110011011010110110000;
   assign mem[202495:202464] = 32'b00000011101000101010000100101000;
   assign mem[202527:202496] = 32'b00000001001110010001111000111100;
   assign mem[202559:202528] = 32'b00000010000101100101000110100100;
   assign mem[202591:202560] = 32'b00001010100011110101001010100000;
   assign mem[202623:202592] = 32'b11101101000010011100011001000000;
   assign mem[202655:202624] = 32'b11111111111110000110100110110101;
   assign mem[202687:202656] = 32'b11111010010111111101110110001000;
   assign mem[202719:202688] = 32'b11100101101000010100011010100000;
   assign mem[202751:202720] = 32'b00000000101110100100110000100000;
   assign mem[202783:202752] = 32'b11111101111101001100110100010100;
   assign mem[202815:202784] = 32'b11110111111000011000011011000000;
   assign mem[202847:202816] = 32'b00000100110001001100001001011000;
   assign mem[202879:202848] = 32'b00000101110100110001110100010000;
   assign mem[202911:202880] = 32'b00000100011101001001100011111000;
   assign mem[202943:202912] = 32'b11110001111011110000111011000000;
   assign mem[202975:202944] = 32'b11111010001001000011110000110000;
   assign mem[203007:202976] = 32'b11111110000100111111101001010110;
   assign mem[203039:203008] = 32'b11111111111100100101010100111110;
   assign mem[203071:203040] = 32'b11110100011010101101011011110000;
   assign mem[203103:203072] = 32'b00000110100000011001101000011000;
   assign mem[203135:203104] = 32'b00000010001110101000010101110000;
   assign mem[203167:203136] = 32'b11111101101010100111000100111100;
   assign mem[203199:203168] = 32'b11111110100110111110011011000100;
   assign mem[203231:203200] = 32'b00000011000001011100100010101000;
   assign mem[203263:203232] = 32'b11110111001110010111111110100000;
   assign mem[203295:203264] = 32'b11111111110011000101010110110010;
   assign mem[203327:203296] = 32'b00000001001001100010000010000110;
   assign mem[203359:203328] = 32'b00000010000110110011010010101100;
   assign mem[203391:203360] = 32'b11110010011101100101000011000000;
   assign mem[203423:203392] = 32'b11111011010000001100011101110000;
   assign mem[203455:203424] = 32'b00000011100010000101110011101100;
   assign mem[203487:203456] = 32'b00000100100001101110110101101000;
   assign mem[203519:203488] = 32'b00000100010111010001111011010000;
   assign mem[203551:203520] = 32'b11110111101010011101010011100000;
   assign mem[203583:203552] = 32'b11111110100111011011111001001000;
   assign mem[203615:203584] = 32'b11111010010110011011111010111000;
   assign mem[203647:203616] = 32'b11101110100011110101001101100000;
   assign mem[203679:203648] = 32'b00000010111100100011011010111100;
   assign mem[203711:203680] = 32'b00000001001110000111010011110110;
   assign mem[203743:203712] = 32'b00000011110100101001000101010000;
   assign mem[203775:203744] = 32'b00000100110010011011110011000000;
   assign mem[203807:203776] = 32'b00000101101111101001010000101000;
   assign mem[203839:203808] = 32'b11110011100010010111111100110000;
   assign mem[203871:203840] = 32'b11110100010111110101110000010000;
   assign mem[203903:203872] = 32'b00001001000111110011001011110000;
   assign mem[203935:203904] = 32'b11111101011010100110000110111000;
   assign mem[203967:203936] = 32'b11111000010111111001100000101000;
   assign mem[203999:203968] = 32'b00001000010010001010000011110000;
   assign mem[204031:204000] = 32'b00000000001101000001000110010001;
   assign mem[204063:204032] = 32'b00000010110101111100011011111100;
   assign mem[204095:204064] = 32'b00000101000101011111010011100000;
   assign mem[204127:204096] = 32'b00000100011100010110110001110000;
   assign mem[204159:204128] = 32'b11110001000001001111011011110000;
   assign mem[204191:204160] = 32'b00000101001000101110010011100000;
   assign mem[204223:204192] = 32'b00000110010110001000100011111000;
   assign mem[204255:204224] = 32'b00000101010111100000001111001000;
   assign mem[204287:204256] = 32'b11110100000110100111000000000000;
   assign mem[204319:204288] = 32'b00001001110000010000000001100000;
   assign mem[204351:204320] = 32'b11101111100110100000011111000000;
   assign mem[204383:204352] = 32'b11110111101010100110011111000000;
   assign mem[204415:204384] = 32'b11111000001001000001111100001000;
   assign mem[204447:204416] = 32'b11111100001100110000100010100100;
   assign mem[204479:204448] = 32'b11110100001111101101111100010000;
   assign mem[204511:204480] = 32'b00000010010111001010100101001100;
   assign mem[204543:204512] = 32'b00000001011111110100101100011110;
   assign mem[204575:204544] = 32'b00001000001001001111000010000000;
   assign mem[204607:204576] = 32'b11111100110101101101101100000100;
   assign mem[204639:204608] = 32'b00000100101100110110100100100000;
   assign mem[204671:204640] = 32'b11110110001000100110101101010000;
   assign mem[204703:204672] = 32'b11110110001110010001001001000000;
   assign mem[204735:204704] = 32'b11111111100100101110010111001000;
   assign mem[204767:204736] = 32'b11111011111001111011000000011000;
   assign mem[204799:204768] = 32'b11111011010101101011100010101000;
   assign mem[204831:204800] = 32'b11110101001000000011100000100000;
   assign mem[204863:204832] = 32'b00000100110110000001001110000000;
   assign mem[204895:204864] = 32'b11111110100111111010000100001110;
   assign mem[204927:204896] = 32'b00000000010011011000000100110000;
   assign mem[204959:204928] = 32'b11111000010111010001111010101000;
   assign mem[204991:204960] = 32'b00000010110010010101101000010000;
   assign mem[205023:204992] = 32'b11111001010101100100011100101000;
   assign mem[205055:205024] = 32'b11111100111100111101111001010000;
   assign mem[205087:205056] = 32'b00000011111001001111011111010000;
   assign mem[205119:205088] = 32'b00000001010110010011110001011000;
   assign mem[205151:205120] = 32'b11110110000000010110010101010000;
   assign mem[205183:205152] = 32'b11110110110110010101100111000000;
   assign mem[205215:205184] = 32'b00000010011011001111110100101000;
   assign mem[205247:205216] = 32'b00000110110000011011100101110000;
   assign mem[205279:205248] = 32'b11111101110010111101010010111000;
   assign mem[205311:205280] = 32'b00000101101101000100111011010000;
   assign mem[205343:205312] = 32'b11111101110111101111011000100000;
   assign mem[205375:205344] = 32'b00000011101110011010110110010000;
   assign mem[205407:205376] = 32'b00000000010011101101000100011110;
   assign mem[205439:205408] = 32'b11111111000011001000000011100011;
   assign mem[205471:205440] = 32'b11111111101100010011011011010001;
   assign mem[205503:205472] = 32'b11110101110010110110011010010000;
   assign mem[205535:205504] = 32'b11110011100000010100101111110000;
   assign mem[205567:205536] = 32'b11110010011110100010111001100000;
   assign mem[205599:205568] = 32'b00000100100100101000011101001000;
   assign mem[205631:205600] = 32'b11111000110010111011010001100000;
   assign mem[205663:205632] = 32'b00000011001110001101010100011100;
   assign mem[205695:205664] = 32'b11111000011010001001001011010000;
   assign mem[205727:205696] = 32'b00001011110111001101110000100000;
   assign mem[205759:205728] = 32'b00000011010111101111100000010100;
   assign mem[205791:205760] = 32'b11110100101011110011010000110000;
   assign mem[205823:205792] = 32'b11111110110001000100001101010100;
   assign mem[205855:205824] = 32'b00000001111010101010001110111000;
   assign mem[205887:205856] = 32'b00000000000011001001100000100100;
   assign mem[205919:205888] = 32'b11111011001110111101101000111000;
   assign mem[205951:205920] = 32'b11111101110110111100000000100000;
   assign mem[205983:205952] = 32'b11101100110001000010100111000000;
   assign mem[206015:205984] = 32'b00000110011101010011111001001000;
   assign mem[206047:206016] = 32'b00000100111010000001110001001000;
   assign mem[206079:206048] = 32'b11110010011001101001110010100000;
   assign mem[206111:206080] = 32'b11111000111110000111011110111000;
   assign mem[206143:206112] = 32'b00000101110000111100101011110000;
   assign mem[206175:206144] = 32'b00001000010011010111111011100000;
   assign mem[206207:206176] = 32'b00000101010110011100111111110000;
   assign mem[206239:206208] = 32'b11110011000000000100110011100000;
   assign mem[206271:206240] = 32'b00000010010100000110101000110000;
   assign mem[206303:206272] = 32'b11110101110100111011100101100000;
   assign mem[206335:206304] = 32'b00000100000001100001010001010000;
   assign mem[206367:206336] = 32'b00000010000000101110110111101000;
   assign mem[206399:206368] = 32'b11111100000001000111010111011000;
   assign mem[206431:206400] = 32'b00000011111100100111011111110100;
   assign mem[206463:206432] = 32'b00000101001011110110011000101000;
   assign mem[206495:206464] = 32'b11110101101010011101001100010000;
   assign mem[206527:206496] = 32'b11110110000111000101101000010000;
   assign mem[206559:206528] = 32'b11111101101101000110011101000000;
   assign mem[206591:206560] = 32'b11111010100110111111101100011000;
   assign mem[206623:206592] = 32'b00001000011100011101011011000000;
   assign mem[206655:206624] = 32'b11110111100100111111110100010000;
   assign mem[206687:206656] = 32'b00000111000110110101110010111000;
   assign mem[206719:206688] = 32'b00000100000101001111111010000000;
   assign mem[206751:206720] = 32'b11111101011111110010000101010100;
   assign mem[206783:206752] = 32'b00000011101111010011000000101000;
   assign mem[206815:206784] = 32'b00000000111101101111011111101110;
   assign mem[206847:206816] = 32'b00000010101011100011010110011000;
   assign mem[206879:206848] = 32'b11111000100001100110000101101000;
   assign mem[206911:206880] = 32'b11111111101111101111100010111001;
   assign mem[206943:206912] = 32'b00000001101001101101110110011010;
   assign mem[206975:206944] = 32'b11110111110010101010011000110000;
   assign mem[207007:206976] = 32'b11111101110011100001010010001100;
   assign mem[207039:207008] = 32'b00000011010011110010000010011000;
   assign mem[207071:207040] = 32'b11111101111000010101110000111100;
   assign mem[207103:207072] = 32'b00000100111110000110001100000000;
   assign mem[207135:207104] = 32'b00000000111010111111011001111101;
   assign mem[207167:207136] = 32'b00000111000100000011011111110000;
   assign mem[207199:207168] = 32'b11110011010011111001010011110000;
   assign mem[207231:207200] = 32'b11110110110101010110010001100000;
   assign mem[207263:207232] = 32'b00000110011110110111010101001000;
   assign mem[207295:207264] = 32'b00000001111000111100101011111100;
   assign mem[207327:207296] = 32'b11110011111011110011010001110000;
   assign mem[207359:207328] = 32'b00000001101011011101110111001100;
   assign mem[207391:207360] = 32'b11111010110111110001110110110000;
   assign mem[207423:207392] = 32'b11111001001011011110000011010000;
   assign mem[207455:207424] = 32'b00001000101000001001111011000000;
   assign mem[207487:207456] = 32'b00000111010010100010110101100000;
   assign mem[207519:207488] = 32'b11111011001011011110001111101000;
   assign mem[207551:207520] = 32'b00000001111100010011010010001010;
   assign mem[207583:207552] = 32'b11110010000101111001010011010000;
   assign mem[207615:207584] = 32'b00000111100110011010101001011000;
   assign mem[207647:207616] = 32'b00000001110101110000110100100100;
   assign mem[207679:207648] = 32'b11110011100110000010010100010000;
   assign mem[207711:207680] = 32'b00000110001000010000000011111000;
   assign mem[207743:207712] = 32'b11110110100110111011011001100000;
   assign mem[207775:207744] = 32'b11111011110110101100100001000000;
   assign mem[207807:207776] = 32'b11110110100101100111011010000000;
   assign mem[207839:207808] = 32'b00000010110101001101101111000100;
   assign mem[207871:207840] = 32'b11111111011111000011010011001100;
   assign mem[207903:207872] = 32'b00001001101101110111000111100000;
   assign mem[207935:207904] = 32'b00000011101011010101001011111100;
   assign mem[207967:207936] = 32'b00000011010111110111110011001100;
   assign mem[207999:207968] = 32'b00000010011000110001101111110000;
   assign mem[208031:208000] = 32'b11111111110000011111000000111010;
   assign mem[208063:208032] = 32'b00000010100111011001000101100000;
   assign mem[208095:208064] = 32'b00000101001010111101101111110000;
   assign mem[208127:208096] = 32'b11111110100010000001100100000010;
   assign mem[208159:208128] = 32'b00000111011000011010111100001000;
   assign mem[208191:208160] = 32'b11110010001100101001011101110000;
   assign mem[208223:208192] = 32'b00000010000101111010111000000000;
   assign mem[208255:208224] = 32'b00000101001111001100100101011000;
   assign mem[208287:208256] = 32'b11111110000110100001100010110010;
   assign mem[208319:208288] = 32'b11111011111110010010010110110000;
   assign mem[208351:208320] = 32'b11111111011100111101010000101110;
   assign mem[208383:208352] = 32'b11111001001101101100001110001000;
   assign mem[208415:208384] = 32'b11111101110110101111100100001100;
   assign mem[208447:208416] = 32'b11111001100111100100011100111000;
   assign mem[208479:208448] = 32'b00000011100100001111110011000000;
   assign mem[208511:208480] = 32'b11111111101111010110100010000111;
   assign mem[208543:208512] = 32'b00000010100010010011001111010100;
   assign mem[208575:208544] = 32'b11111001011101110100010001111000;
   assign mem[208607:208576] = 32'b00000100010110001011101111011000;
   assign mem[208639:208608] = 32'b00000110001001101101100001100000;
   assign mem[208671:208640] = 32'b11111100010110011000101100001000;
   assign mem[208703:208672] = 32'b11111101100010101000011000000100;
   assign mem[208735:208704] = 32'b00001010001101010100010101100000;
   assign mem[208767:208736] = 32'b11111001101111110111011111111000;
   assign mem[208799:208768] = 32'b11110010010001001100011001010000;
   assign mem[208831:208800] = 32'b00000010000111110110111001110100;
   assign mem[208863:208832] = 32'b11111010010111111110010111100000;
   assign mem[208895:208864] = 32'b11101111111000101011010000000000;
   assign mem[208927:208896] = 32'b00001000011110110110010011010000;
   assign mem[208959:208928] = 32'b11111110010101101011101000000100;
   assign mem[208991:208960] = 32'b11110100111110100111010100100000;
   assign mem[209023:208992] = 32'b11110100111110100000000000010000;
   assign mem[209055:209024] = 32'b00000110010001001101110101010000;
   assign mem[209087:209056] = 32'b00001001100010111011001000110000;
   assign mem[209119:209088] = 32'b11111000011100011100000010011000;
   assign mem[209151:209120] = 32'b00000100000101001110100110100000;
   assign mem[209183:209152] = 32'b11110001100000100001011000000000;
   assign mem[209215:209184] = 32'b00000001111000000001001100010100;
   assign mem[209247:209216] = 32'b00000000010100111010010000010110;
   assign mem[209279:209248] = 32'b11110111001101000010011111110000;
   assign mem[209311:209280] = 32'b00000001011000010110101000111110;
   assign mem[209343:209312] = 32'b11111001000111001101100101011000;
   assign mem[209375:209344] = 32'b11111100011101111111110101010100;
   assign mem[209407:209376] = 32'b11110011010011011011011110100000;
   assign mem[209439:209408] = 32'b00000011001010100100010011001000;
   assign mem[209471:209440] = 32'b00000001101101101110010001100100;
   assign mem[209503:209472] = 32'b00000100101100100101101101101000;
   assign mem[209535:209504] = 32'b11111000001010010001000110011000;
   assign mem[209567:209536] = 32'b00000101101110001111000111000000;
   assign mem[209599:209568] = 32'b00000110100101010000010011011000;
   assign mem[209631:209600] = 32'b00000100101010000000000011011000;
   assign mem[209663:209632] = 32'b11111101011000110100101001101100;
   assign mem[209695:209664] = 32'b11111101111110100101111101001000;
   assign mem[209727:209696] = 32'b11110011001110001100100010010000;
   assign mem[209759:209728] = 32'b11111111000110111001011001100011;
   assign mem[209791:209760] = 32'b11111111100111101011011110100000;
   assign mem[209823:209792] = 32'b00000101010011010100011100111000;
   assign mem[209855:209824] = 32'b11111111011011111001100111101111;
   assign mem[209887:209856] = 32'b00000000000110101110010100011010;
   assign mem[209919:209888] = 32'b00000011001110000101100011111100;
   assign mem[209951:209920] = 32'b11111010110100101100010000100000;
   assign mem[209983:209952] = 32'b11111010101110000110000100100000;
   assign mem[210015:209984] = 32'b00000100101110000100011010111000;
   assign mem[210047:210016] = 32'b00000101111010101110101000000000;
   assign mem[210079:210048] = 32'b11111111010010110101011011000000;
   assign mem[210111:210080] = 32'b00000010110110101111011010101100;
   assign mem[210143:210112] = 32'b11101111010000111111100011100000;
   assign mem[210175:210144] = 32'b00000101110010100011011101100000;
   assign mem[210207:210176] = 32'b11111001001011001001000010111000;
   assign mem[210239:210208] = 32'b11111001001000001100100110100000;
   assign mem[210271:210240] = 32'b11111110110010101100001100111000;
   assign mem[210303:210272] = 32'b11111110100011010101100001010010;
   assign mem[210335:210304] = 32'b11110001101010010100010101000000;
   assign mem[210367:210336] = 32'b11111010000100110010101100010000;
   assign mem[210399:210368] = 32'b00000000100111100101001100001110;
   assign mem[210431:210400] = 32'b11111010101100001111010110010000;
   assign mem[210463:210432] = 32'b00000100110000101101001001110000;
   assign mem[210495:210464] = 32'b00000000000100101111011000001110;
   assign mem[210527:210496] = 32'b00000100010000001000001110001000;
   assign mem[210559:210528] = 32'b00000010110101110111011000111100;
   assign mem[210591:210560] = 32'b11111000110011001000010101011000;
   assign mem[210623:210592] = 32'b11110111110000101001101100100000;
   assign mem[210655:210624] = 32'b00000011010001011001010111001100;
   assign mem[210687:210656] = 32'b00000110101000011111011011000000;
   assign mem[210719:210688] = 32'b11111000011111100110001011100000;
   assign mem[210751:210720] = 32'b11111001000100000100101000000000;
   assign mem[210783:210752] = 32'b11110100010110101111101111010000;
   assign mem[210815:210784] = 32'b00000010000000110011001011100000;
   assign mem[210847:210816] = 32'b00000011100000000101100110100100;
   assign mem[210879:210848] = 32'b11111000000100100001110011110000;
   assign mem[210911:210880] = 32'b00000100111010110010001010001000;
   assign mem[210943:210912] = 32'b11111000100110100000011101100000;
   assign mem[210975:210944] = 32'b00001100010000111100101100010000;
   assign mem[211007:210976] = 32'b00000011100001001010011001100000;
   assign mem[211039:211008] = 32'b00000101101010100010001101110000;
   assign mem[211071:211040] = 32'b11111000101111101010101000101000;
   assign mem[211103:211072] = 32'b11111011000101101100101110011000;
   assign mem[211135:211104] = 32'b11111011110001011011100000110000;
   assign mem[211167:211136] = 32'b11111110111101000010100101010110;
   assign mem[211199:211168] = 32'b11110100110001011011000100010000;
   assign mem[211231:211200] = 32'b00000100111101000001100010101000;
   assign mem[211263:211232] = 32'b00000001111110001001101111101110;
   assign mem[211295:211264] = 32'b11110001100100000101100001100000;
   assign mem[211327:211296] = 32'b11111001001010100001101001001000;
   assign mem[211359:211328] = 32'b00000001100111010111111111101010;
   assign mem[211391:211360] = 32'b11111111100100011110101100111001;
   assign mem[211423:211392] = 32'b00000010100011000001011011101000;
   assign mem[211455:211424] = 32'b00001000100111111111011001100000;
   assign mem[211487:211456] = 32'b11111111111100001000110000011000;
   assign mem[211519:211488] = 32'b00000100101001010000100001011000;
   assign mem[211551:211520] = 32'b00000011010011110101010001010100;
   assign mem[211583:211552] = 32'b11111101110111101011001100110100;
   assign mem[211615:211584] = 32'b00001001001110010110000001000000;
   assign mem[211647:211616] = 32'b00000001010000100110010011011110;
   assign mem[211679:211648] = 32'b00000010011111110010101001111100;
   assign mem[211711:211680] = 32'b11110010001100010000001110110000;
   assign mem[211743:211712] = 32'b11110100000011011101011110110000;
   assign mem[211775:211744] = 32'b00000111100010101110111011101000;
   assign mem[211807:211776] = 32'b11111110110110010111001000010010;
   assign mem[211839:211808] = 32'b11101110001111000111101001000000;
   assign mem[211871:211840] = 32'b00000010011010010011100111111100;
   assign mem[211903:211872] = 32'b00000010011101100011011010110100;
   assign mem[211935:211904] = 32'b11111101000011000100010000000000;
   assign mem[211967:211936] = 32'b11111000010100001101000110000000;
   assign mem[211999:211968] = 32'b00000011010000100000010101000000;
   assign mem[212031:212000] = 32'b11111100001000111111111111011100;
   assign mem[212063:212032] = 32'b00000100001001010010000000001000;
   assign mem[212095:212064] = 32'b11111111001101111011110001001111;
   assign mem[212127:212096] = 32'b11110110100111011101100100000000;
   assign mem[212159:212128] = 32'b00000100110101101101000100001000;
   assign mem[212191:212160] = 32'b00000110011011111100111110001000;
   assign mem[212223:212192] = 32'b11110111010011101111110101010000;
   assign mem[212255:212224] = 32'b11101111110111111101100001000000;
   assign mem[212287:212256] = 32'b11111001100011110110100110110000;
   assign mem[212319:212288] = 32'b00000110110011011010010111111000;
   assign mem[212351:212320] = 32'b11111111000100011110110010110000;
   assign mem[212383:212352] = 32'b00000001111101100110100011000100;
   assign mem[212415:212384] = 32'b11111101011101111100011001100100;
   assign mem[212447:212416] = 32'b00000110010100001101101100011000;
   assign mem[212479:212448] = 32'b00001001000100000111011110000000;
   assign mem[212511:212480] = 32'b00000001011100011001101100100010;
   assign mem[212543:212512] = 32'b11111001001111110011111100011000;
   assign mem[212575:212544] = 32'b11111011101101011011111000100000;
   assign mem[212607:212576] = 32'b11111001111100011100111010111000;
   assign mem[212639:212608] = 32'b11111100011110100101100110101100;
   assign mem[212671:212640] = 32'b00000000001100101011110100010111;
   assign mem[212703:212672] = 32'b00000100011101110111010100101000;
   assign mem[212735:212704] = 32'b11111011101010001011110001100000;
   assign mem[212767:212736] = 32'b00000110001000000100010111101000;
   assign mem[212799:212768] = 32'b00000111010101000101011101000000;
   assign mem[212831:212800] = 32'b00000000000001110001101110011000;
   assign mem[212863:212832] = 32'b00000100110100110001000010000000;
   assign mem[212895:212864] = 32'b11111101011001111000101001010000;
   assign mem[212927:212896] = 32'b00000010001100010000001000011000;
   assign mem[212959:212928] = 32'b11111001110000101000010101111000;
   assign mem[212991:212960] = 32'b11110101101000100000000001100000;
   assign mem[213023:212992] = 32'b00001101010100000010000001010000;
   assign mem[213055:213024] = 32'b11111011101011011010100110000000;
   assign mem[213087:213056] = 32'b11110101010001110001001100010000;
   assign mem[213119:213088] = 32'b00000100001001001011000011000000;
   assign mem[213151:213120] = 32'b11111010000110010011111111001000;
   assign mem[213183:213152] = 32'b00000100000110010111001101111000;
   assign mem[213215:213184] = 32'b11101111101111110000010001000000;
   assign mem[213247:213216] = 32'b00000101001010000111100011100000;
   assign mem[213279:213248] = 32'b11110011101001101000110100110000;
   assign mem[213311:213280] = 32'b11111110101001001000110111110010;
   assign mem[213343:213312] = 32'b00000110001000100010000000000000;
   assign mem[213375:213344] = 32'b11110110100011110001000111010000;
   assign mem[213407:213376] = 32'b11111110101001001001110011101000;
   assign mem[213439:213408] = 32'b00000100001100100111110010001000;
   assign mem[213471:213440] = 32'b00000100001111101000100110110000;
   assign mem[213503:213472] = 32'b11111011011000001100010001000000;
   assign mem[213535:213504] = 32'b00000010110110101110011001100100;
   assign mem[213567:213536] = 32'b11111001100100111111100011111000;
   assign mem[213599:213568] = 32'b00000000011100100010101110011010;
   assign mem[213631:213600] = 32'b00000001000011011001000111111010;
   assign mem[213663:213632] = 32'b11111110101101111100101110000110;
   assign mem[213695:213664] = 32'b11111010010110110011001010111000;
   assign mem[213727:213696] = 32'b11111110100110100001100101111100;
   assign mem[213759:213728] = 32'b11111010110001000100100111100000;
   assign mem[213791:213760] = 32'b11111100111111001111001011100000;
   assign mem[213823:213792] = 32'b00000001111101001101100000010100;
   assign mem[213855:213824] = 32'b00000010000100010010101000001000;
   assign mem[213887:213856] = 32'b11111010001101110001110110111000;
   assign mem[213919:213888] = 32'b11111100101011010000010011100100;
   assign mem[213951:213920] = 32'b11111100101100010011011100011000;
   assign mem[213983:213952] = 32'b00000000011011111010001011111001;
   assign mem[214015:213984] = 32'b00000010100111100111000111100100;
   assign mem[214047:214016] = 32'b00000000111101011100100011110110;
   assign mem[214079:214048] = 32'b00000100100111101100000100010000;
   assign mem[214111:214080] = 32'b11111000100001110110101010001000;
   assign mem[214143:214112] = 32'b11111001101100001111100001000000;
   assign mem[214175:214144] = 32'b00001001100100010001111011000000;
   assign mem[214207:214176] = 32'b00000011100111100110110110110100;
   assign mem[214239:214208] = 32'b11111011110000010010010101101000;
   assign mem[214271:214240] = 32'b11111111101111001111010001010101;
   assign mem[214303:214272] = 32'b11110010001110100101011111110000;
   assign mem[214335:214304] = 32'b00001001111111110100000100000000;
   assign mem[214367:214336] = 32'b00000101101111001010011000100000;
   assign mem[214399:214368] = 32'b11101110010110001111101001000000;
   assign mem[214431:214400] = 32'b00000100111010000110000101011000;
   assign mem[214463:214432] = 32'b00000001000100000101100110011010;
   assign mem[214495:214464] = 32'b11101110000101111011010001100000;
   assign mem[214527:214496] = 32'b00000110101100000010111010010000;
   assign mem[214559:214528] = 32'b00001010001010000000010110000000;
   assign mem[214591:214560] = 32'b11110000010100101001000110010000;
   assign mem[214623:214592] = 32'b00000000011001111100000000011000;
   assign mem[214655:214624] = 32'b00000100011101000110000100100000;
   assign mem[214687:214656] = 32'b11111000101100111111111100101000;
   assign mem[214719:214688] = 32'b11111110100111011111000011000000;
   assign mem[214751:214720] = 32'b11110101101111111001101111100000;
   assign mem[214783:214752] = 32'b11110101000000010001110011100000;
   assign mem[214815:214784] = 32'b00000100111101010100111000011000;
   assign mem[214847:214816] = 32'b00000100000100001101101010001000;
   assign mem[214879:214848] = 32'b00000100110011011110101100110000;
   assign mem[214911:214880] = 32'b00000001111010101010000010110010;
   assign mem[214943:214912] = 32'b11110001100111111000111001010000;
   assign mem[214975:214944] = 32'b00000011000111010010110111010000;
   assign mem[215007:214976] = 32'b00000001001001011010110001101010;
   assign mem[215039:215008] = 32'b11111111110010000000110010001001;
   assign mem[215071:215040] = 32'b00000101000010010100110000000000;
   assign mem[215103:215072] = 32'b11111100010001101101010111010100;
   assign mem[215135:215104] = 32'b11111111100011011101000110100001;
   assign mem[215167:215136] = 32'b11111011010101110000110011000000;
   assign mem[215199:215168] = 32'b00000001000001100001100101000000;
   assign mem[215231:215200] = 32'b11110001000001110011101000110000;
   assign mem[215263:215232] = 32'b00001001110010111101101001110000;
   assign mem[215295:215264] = 32'b00000001011010100011101110000100;
   assign mem[215327:215296] = 32'b00000011001010110001010110101100;
   assign mem[215359:215328] = 32'b00000011000100111111001110101000;
   assign mem[215391:215360] = 32'b00000101101111100101001000001000;
   assign mem[215423:215392] = 32'b00000011101100110111110100001100;
   assign mem[215455:215424] = 32'b11110101000110011001011001010000;
   assign mem[215487:215456] = 32'b11111011011111100101111111010000;
   assign mem[215519:215488] = 32'b11111101101010100000001100000000;
   assign mem[215551:215520] = 32'b11111000001001100001010111110000;
   assign mem[215583:215552] = 32'b00000011110001110111101011011000;
   assign mem[215615:215584] = 32'b11111111011111011101001110100010;
   assign mem[215647:215616] = 32'b00000011000001110110110000000000;
   assign mem[215679:215648] = 32'b00000100111001100011110110111000;
   assign mem[215711:215680] = 32'b11110010110001101110010001100000;
   assign mem[215743:215712] = 32'b11110111001010011101110000100000;
   assign mem[215775:215744] = 32'b00000011011010010001001011000000;
   assign mem[215807:215776] = 32'b11110100000001001101110011110000;
   assign mem[215839:215808] = 32'b00000101011110000101011010000000;
   assign mem[215871:215840] = 32'b00000000100000100000010001001000;
   assign mem[215903:215872] = 32'b11111100100000001000000111110100;
   assign mem[215935:215904] = 32'b11111011111001111001010111110000;
   assign mem[215967:215936] = 32'b11111110110010101100101011010010;
   assign mem[215999:215968] = 32'b00001000011001111000100100000000;
   assign mem[216031:216000] = 32'b00000100000111000011111001010000;
   assign mem[216063:216032] = 32'b11111010010111011010001110101000;
   assign mem[216095:216064] = 32'b00000111001001000111011110001000;
   assign mem[216127:216096] = 32'b11111000110100010011001000000000;
   assign mem[216159:216128] = 32'b00000000111100100001101110010110;
   assign mem[216191:216160] = 32'b00000010010110110100010001110000;
   assign mem[216223:216192] = 32'b11111100100111110011111100000100;
   assign mem[216255:216224] = 32'b11111000110000101101110100111000;
   assign mem[216287:216256] = 32'b11111101110111110111011010110100;
   assign mem[216319:216288] = 32'b11111110100111001000001001011100;
   assign mem[216351:216320] = 32'b11101001011010000001010001100000;
   assign mem[216383:216352] = 32'b11111110111000110111101000000100;
   assign mem[216415:216384] = 32'b00000011110011011010110110011100;
   assign mem[216447:216416] = 32'b00000111100101011001001110111000;
   assign mem[216479:216448] = 32'b11110100100000110110100011000000;
   assign mem[216511:216480] = 32'b00000011111011100100111001000100;
   assign mem[216543:216512] = 32'b11101101111100010011111100000000;
   assign mem[216575:216544] = 32'b00000010100110110000100010100100;
   assign mem[216607:216576] = 32'b00000010111101110011110101101000;
   assign mem[216639:216608] = 32'b11111110011000000100110100111100;
   assign mem[216671:216640] = 32'b11111000001010010011011001111000;
   assign mem[216703:216672] = 32'b11111101011111101011010110100100;
   assign mem[216735:216704] = 32'b00000111000001111011111011110000;
   assign mem[216767:216736] = 32'b00000111100110111000101010010000;
   assign mem[216799:216768] = 32'b11111010000100000110110011110000;
   assign mem[216831:216800] = 32'b11111011011111010111000001101000;
   assign mem[216863:216832] = 32'b00000110011110000010100100101000;
   assign mem[216895:216864] = 32'b00001000100010001100101000100000;
   assign mem[216927:216896] = 32'b00000001111110100100001001111000;
   assign mem[216959:216928] = 32'b11111110010001010110100100101110;
   assign mem[216991:216960] = 32'b11111000001000001101110100100000;
   assign mem[217023:216992] = 32'b00000000100011110111111110100110;
   assign mem[217055:217024] = 32'b11111001000000001110001100111000;
   assign mem[217087:217056] = 32'b11101111100010111100001110000000;
   assign mem[217119:217088] = 32'b00001001001001101001001110110000;
   assign mem[217151:217120] = 32'b00000001101001101011001101101000;
   assign mem[217183:217152] = 32'b00000100010010001111101110010000;
   assign mem[217215:217184] = 32'b11111100001101010111110100010100;
   assign mem[217247:217216] = 32'b00000100000011000010101101110000;
   assign mem[217279:217248] = 32'b00000010010111101001101101011000;
   assign mem[217311:217280] = 32'b00000010011000101100001000000100;
   assign mem[217343:217312] = 32'b11111010011101101111110110000000;
   assign mem[217375:217344] = 32'b00001000110101110001111111010000;
   assign mem[217407:217376] = 32'b00000100010101011010101000001000;
   assign mem[217439:217408] = 32'b11111001010101100111111110100000;
   assign mem[217471:217440] = 32'b11111011011011010001110001110000;
   assign mem[217503:217472] = 32'b11111100011011111010110000010000;
   assign mem[217535:217504] = 32'b11111101001011100010010100000100;
   assign mem[217567:217536] = 32'b00000100001100110001110011100000;
   assign mem[217599:217568] = 32'b11101110000100100001110011000000;
   assign mem[217631:217600] = 32'b11111101110010110000001001111000;
   assign mem[217663:217632] = 32'b11110111111100110101100001100000;
   assign mem[217695:217664] = 32'b11111100101000100011110101100100;
   assign mem[217727:217696] = 32'b11101101001100010011111111000000;
   assign mem[217759:217728] = 32'b00000110001100111100110011111000;
   assign mem[217791:217760] = 32'b00000001011010000100000111100100;
   assign mem[217823:217792] = 32'b00000000011101011111011000111100;
   assign mem[217855:217824] = 32'b11111001011101100011001101000000;
   assign mem[217887:217856] = 32'b00000011100010000111001010001000;
   assign mem[217919:217888] = 32'b00001001000010111101101010010000;
   assign mem[217951:217920] = 32'b11111101001101001100000111001100;
   assign mem[217983:217952] = 32'b00001000101111110000110111000000;
   assign mem[218015:217984] = 32'b00000101001010101100110010001000;
   assign mem[218047:218016] = 32'b00000011001101011000100101000100;
   assign mem[218079:218048] = 32'b11110000100111100011001000110000;
   assign mem[218111:218080] = 32'b11111110000100101000110010101110;
   assign mem[218143:218112] = 32'b11111001001111001010101101001000;
   assign mem[218175:218144] = 32'b00001001001101000100001101110000;
   assign mem[218207:218176] = 32'b11111101001111000000100000100000;
   assign mem[218239:218208] = 32'b11111001000010101011101111010000;
   assign mem[218271:218240] = 32'b11110111001100001011000111100000;
   assign mem[218303:218272] = 32'b00000100001111111000111110001000;
   assign mem[218335:218304] = 32'b00000000011101110011001111010011;
   assign mem[218367:218336] = 32'b00000011100011111100010011111100;
   assign mem[218399:218368] = 32'b11111100001101110110010011001100;
   assign mem[218431:218400] = 32'b11111111010100010011000010101011;
   assign mem[218463:218432] = 32'b11101001011110110110100010100000;
   assign mem[218495:218464] = 32'b00000001000110111100011110100010;
   assign mem[218527:218496] = 32'b00000010011000001011011100001100;
   assign mem[218559:218528] = 32'b11111101111010011101011101111000;
   assign mem[218591:218560] = 32'b11111010010001001111001001110000;
   assign mem[218623:218592] = 32'b00000010011000011110100000010100;
   assign mem[218655:218624] = 32'b11111011000001010001110000000000;
   assign mem[218687:218656] = 32'b00000001001100110100011000100100;
   assign mem[218719:218688] = 32'b00000011111100001010010100110000;
   assign mem[218751:218720] = 32'b11111110001100000010011010001100;
   assign mem[218783:218752] = 32'b00000100001000110101110001111000;
   assign mem[218815:218784] = 32'b00001000111001101110000000110000;
   assign mem[218847:218816] = 32'b11111110111100011110001101101000;
   assign mem[218879:218848] = 32'b00000010101101011110101001101100;
   assign mem[218911:218880] = 32'b00000000010100001011111010100010;
   assign mem[218943:218912] = 32'b11111000100100101100001001111000;
   assign mem[218975:218944] = 32'b11110111111101100101110010100000;
   assign mem[219007:218976] = 32'b11101111101101010101111111100000;
   assign mem[219039:219008] = 32'b00001001111100011001010011000000;
   assign mem[219071:219040] = 32'b00000010000010111110111001110100;
   assign mem[219103:219072] = 32'b11111001010111010001100100111000;
   assign mem[219135:219104] = 32'b11110011110010010001010100010000;
   assign mem[219167:219136] = 32'b00000011011111000101110010111000;
   assign mem[219199:219168] = 32'b00001001101011011101110000110000;
   assign mem[219231:219200] = 32'b00000010100110111100001010111100;
   assign mem[219263:219232] = 32'b11111011101110000110110011000000;
   assign mem[219295:219264] = 32'b00000101000001001001110011111000;
   assign mem[219327:219296] = 32'b11111110110011111011000101011010;
   assign mem[219359:219328] = 32'b00000011000011011100010101101000;
   assign mem[219391:219360] = 32'b11111100111101110010110001101000;
   assign mem[219423:219392] = 32'b00000000011000100010001100111001;
   assign mem[219455:219424] = 32'b00000100010001010100101010001000;
   assign mem[219487:219456] = 32'b11111100111111000011110110101000;
   assign mem[219519:219488] = 32'b00000000010010010001011001110100;
   assign mem[219551:219520] = 32'b00000000001101111100010111011111;
   assign mem[219583:219552] = 32'b11111010100101011010000001110000;
   assign mem[219615:219584] = 32'b11111010001010101000011101010000;
   assign mem[219647:219616] = 32'b11111010001110100000011100101000;
   assign mem[219679:219648] = 32'b11111100111100001101110111111000;
   assign mem[219711:219680] = 32'b00000011000011101100101000101100;
   assign mem[219743:219712] = 32'b00000001101100000110000110110000;
   assign mem[219775:219744] = 32'b00000110011110110110010111100000;
   assign mem[219807:219776] = 32'b00000011010111010111011101100000;
   assign mem[219839:219808] = 32'b00000001010101111001001011101110;
   assign mem[219871:219840] = 32'b11111101110001101010101100100100;
   assign mem[219903:219872] = 32'b11111011111010100000010010000000;
   assign mem[219935:219904] = 32'b11111111010101111110110110001101;
   assign mem[219967:219936] = 32'b00000001001001111010011001000100;
   assign mem[219999:219968] = 32'b00000010011001100011011000000100;
   assign mem[220031:220000] = 32'b00000001011110111100001011101010;
   assign mem[220063:220032] = 32'b11111110101011011001111101000000;
   assign mem[220095:220064] = 32'b11111111101000001101110110010111;
   assign mem[220127:220096] = 32'b00000010010101100011011110100000;
   assign mem[220159:220128] = 32'b00000001010110111001000000111100;
   assign mem[220191:220160] = 32'b11110011101101011010011100100000;
   assign mem[220223:220192] = 32'b11111101111000110110101010101000;
   assign mem[220255:220224] = 32'b11110011100100010010110010000000;
   assign mem[220287:220256] = 32'b11110101011111000101011001010000;
   assign mem[220319:220288] = 32'b11111100111000101001100010011000;
   assign mem[220351:220320] = 32'b11111101001100110101101100010100;
   assign mem[220383:220352] = 32'b11111001011001100001101010101000;
   assign mem[220415:220384] = 32'b00010001000010011000000101000000;
   assign mem[220447:220416] = 32'b00000100010111010101101110101000;
   assign mem[220479:220448] = 32'b11111110011111011100011001000110;
   assign mem[220511:220480] = 32'b00001000000011101111000110110000;
   assign mem[220543:220512] = 32'b11110100111111101101000101000000;
   assign mem[220575:220544] = 32'b00000001111100101110101111100100;
   assign mem[220607:220576] = 32'b11101111101110000110000111000000;
   assign mem[220639:220608] = 32'b00000101001111110011001011011000;
   assign mem[220671:220640] = 32'b11111001111101100110100001100000;
   assign mem[220703:220672] = 32'b00000101111100111110000011010000;
   assign mem[220735:220704] = 32'b11111111011000010000010010010111;
   assign mem[220767:220736] = 32'b11111110100111000100011100110110;
   assign mem[220799:220768] = 32'b00000100110000011100000010000000;
   assign mem[220831:220800] = 32'b00000011001000100110110010010000;
   assign mem[220863:220832] = 32'b00000001010110101110101110110000;
   assign mem[220895:220864] = 32'b00000000101101101100011111100000;
   assign mem[220927:220896] = 32'b11110111011101000000000011010000;
   assign mem[220959:220928] = 32'b00000000001111101011111011000110;
   assign mem[220991:220960] = 32'b11111010101000100110011000000000;
   assign mem[221023:220992] = 32'b00000111100100100010000011100000;
   assign mem[221055:221024] = 32'b11111110000011000100101100011100;
   assign mem[221087:221056] = 32'b00000111010111101111010001101000;
   assign mem[221119:221088] = 32'b00000100111111001100010001001000;
   assign mem[221151:221120] = 32'b11111111111110010110111010001011;
   assign mem[221183:221152] = 32'b11111101000011100111110111000000;
   assign mem[221215:221184] = 32'b00000001111010101001110111100010;
   assign mem[221247:221216] = 32'b11111111100000101110001011000011;
   assign mem[221279:221248] = 32'b00000000100001111101110101100111;
   assign mem[221311:221280] = 32'b11111111100100011110110011111001;
   assign mem[221343:221312] = 32'b00000010001101100101000100001100;
   assign mem[221375:221344] = 32'b11111100001111011000010011000100;
   assign mem[221407:221376] = 32'b11111110110000101000101110101010;
   assign mem[221439:221408] = 32'b11111010111000000011110011111000;
   assign mem[221471:221440] = 32'b11110111111011011100100010000000;
   assign mem[221503:221472] = 32'b11110110111101010110010101000000;
   assign mem[221535:221504] = 32'b11111111001011000110000111011101;
   assign mem[221567:221536] = 32'b11111111010000101011110101110100;
   assign mem[221599:221568] = 32'b00000100000001110110110111110000;
   assign mem[221631:221600] = 32'b00000110101111011100000101000000;
   assign mem[221663:221632] = 32'b11111010010011001111101101011000;
   assign mem[221695:221664] = 32'b11111101100110010001010011011000;
   assign mem[221727:221696] = 32'b00000101000000101001000000111000;
   assign mem[221759:221728] = 32'b11111110001100100111111111001110;
   assign mem[221791:221760] = 32'b11111001001101010110011110001000;
   assign mem[221823:221792] = 32'b11111110000010011001101111011100;
   assign mem[221855:221824] = 32'b00000000100111101111110100011010;
   assign mem[221887:221856] = 32'b11111101010001001011001000110100;
   assign mem[221919:221888] = 32'b00000111001001010011111010000000;
   assign mem[221951:221920] = 32'b11111011100100100100100111001000;
   assign mem[221983:221952] = 32'b11110100111011011000011110100000;
   assign mem[222015:221984] = 32'b00000010001101010001101110010100;
   assign mem[222047:222016] = 32'b00001001110010110110100110000000;
   assign mem[222079:222048] = 32'b00000001011101100001101100001100;
   assign mem[222111:222080] = 32'b11111001100011101110000010101000;
   assign mem[222143:222112] = 32'b11110111001000101101101100010000;
   assign mem[222175:222144] = 32'b11111110001100010000110111101100;
   assign mem[222207:222176] = 32'b11111110111000111010100110010110;
   assign mem[222239:222208] = 32'b00000100100011000001110110101000;
   assign mem[222271:222240] = 32'b00000111110001011111000101011000;
   assign mem[222303:222272] = 32'b11110001000001100101110000110000;
   assign mem[222335:222304] = 32'b00000001110110100101010001011100;
   assign mem[222367:222336] = 32'b11111111000011110010110010011101;
   assign mem[222399:222368] = 32'b00000111001111010011101100000000;
   assign mem[222431:222400] = 32'b11111111001001010000000100110011;
   assign mem[222463:222432] = 32'b00000100101110010100100000010000;
   assign mem[222495:222464] = 32'b00000000001001110010001000001010;
   assign mem[222527:222496] = 32'b11111100110001110110000000110000;
   assign mem[222559:222528] = 32'b00000010110010011011101011011000;
   assign mem[222591:222560] = 32'b11111110000000100101010001001010;
   assign mem[222623:222592] = 32'b00000101010011001100100101010000;
   assign mem[222655:222624] = 32'b11111100101000100111001011000000;
   assign mem[222687:222656] = 32'b00000010011000011001000000000100;
   assign mem[222719:222688] = 32'b00000100111100111110110000001000;
   assign mem[222751:222720] = 32'b00000000101001100001000110010111;
   assign mem[222783:222752] = 32'b11111110111101111001001100000000;
   assign mem[222815:222784] = 32'b11111101101010100010100100001000;
   assign mem[222847:222816] = 32'b11111110011101110100011001100010;
   assign mem[222879:222848] = 32'b00000001111001101000110010010010;
   assign mem[222911:222880] = 32'b00000000110000110001001010000011;
   assign mem[222943:222912] = 32'b11111101101001101011001000010100;
   assign mem[222975:222944] = 32'b00000110010001001001100101010000;
   assign mem[223007:222976] = 32'b00000000011100111101100101010001;
   assign mem[223039:223008] = 32'b00000010100100010010001100101100;
   assign mem[223071:223040] = 32'b11110011111001011011110001110000;
   assign mem[223103:223072] = 32'b00000001011010101001110110110110;
   assign mem[223135:223104] = 32'b11111100100011001011101011111100;
   assign mem[223167:223136] = 32'b11111101001111001000000011100000;
   assign mem[223199:223168] = 32'b00000100010010111100101011110000;
   assign mem[223231:223200] = 32'b00000011001000001110011001101100;
   assign mem[223263:223232] = 32'b11111111010110111001010100011010;
   assign mem[223295:223264] = 32'b00000000000000111011001000001000;
   assign mem[223327:223296] = 32'b00000011001011000110110110111100;
   assign mem[223359:223328] = 32'b00000111110110100100001000011000;
   assign mem[223391:223360] = 32'b00000011011010011100110000011000;
   assign mem[223423:223392] = 32'b11111001001111001101010100111000;
   assign mem[223455:223424] = 32'b00001000011001000011101000010000;
   assign mem[223487:223456] = 32'b11111111010010111010110001110001;
   assign mem[223519:223488] = 32'b11111100010110001000101000111100;
   assign mem[223551:223520] = 32'b11111101010011110011101111000100;
   assign mem[223583:223552] = 32'b11111110011110010100011101110010;
   assign mem[223615:223584] = 32'b11111110010101100110000100111000;
   assign mem[223647:223616] = 32'b11111101100101011100010011100000;
   assign mem[223679:223648] = 32'b11110110111001111100001101110000;
   assign mem[223711:223680] = 32'b00000101001110000101100110010000;
   assign mem[223743:223712] = 32'b11111110011111100101010110000100;
   assign mem[223775:223744] = 32'b00000111111010110010110100101000;
   assign mem[223807:223776] = 32'b11111111000100000100101011001101;
   assign mem[223839:223808] = 32'b00000111100101110101001011000000;
   assign mem[223871:223840] = 32'b11111001111001111100110110011000;
   assign mem[223903:223872] = 32'b00000000001110101101101011111100;
   assign mem[223935:223904] = 32'b00000001000010001110101010110000;
   assign mem[223967:223936] = 32'b11111100111000010111110010001000;
   assign mem[223999:223968] = 32'b11110011010101100101001101100000;
   assign mem[224031:224000] = 32'b00000011110000001001100011100000;
   assign mem[224063:224032] = 32'b11111100101011101010000001101100;
   assign mem[224095:224064] = 32'b00001010001000110100100100010000;
   assign mem[224127:224096] = 32'b00000001010000001011001110111000;
   assign mem[224159:224128] = 32'b00000000101011100111111100110100;
   assign mem[224191:224160] = 32'b11111110110111000111111101100000;
   assign mem[224223:224192] = 32'b11111100011100110100011100010000;
   assign mem[224255:224224] = 32'b11111101000011111011111011011100;
   assign mem[224287:224256] = 32'b00000001110011110011111010001100;
   assign mem[224319:224288] = 32'b11110110001000010001011100010000;
   assign mem[224351:224320] = 32'b00000010011001011011000100010100;
   assign mem[224383:224352] = 32'b11110011101111011101010110100000;
   assign mem[224415:224384] = 32'b11111111011111010000110001011001;
   assign mem[224447:224416] = 32'b11110011000001101110100010010000;
   assign mem[224479:224448] = 32'b00000100010010101111001001010000;
   assign mem[224511:224480] = 32'b11111001001000010101010111101000;
   assign mem[224543:224512] = 32'b00000100010010011100000111100000;
   assign mem[224575:224544] = 32'b00000011011000111001001101111000;
   assign mem[224607:224576] = 32'b11111110110011000011010000111010;
   assign mem[224639:224608] = 32'b00000100000001010001100011010000;
   assign mem[224671:224640] = 32'b00000100001111010110010001011000;
   assign mem[224703:224672] = 32'b11111001110001001111101010000000;
   assign mem[224735:224704] = 32'b11111100111011010001000101100100;
   assign mem[224767:224736] = 32'b11110011100101000001101110000000;
   assign mem[224799:224768] = 32'b00000000001001101000100000110011;
   assign mem[224831:224800] = 32'b00000001001111110101010001010100;
   assign mem[224863:224832] = 32'b00000100101110100010010001001000;
   assign mem[224895:224864] = 32'b11111111001010110100110000001110;
   assign mem[224927:224896] = 32'b11111111000110000101011100010011;
   assign mem[224959:224928] = 32'b11111111100000111100110101110111;
   assign mem[224991:224960] = 32'b00000010101010110100110000111100;
   assign mem[225023:224992] = 32'b11101111010101000111100011000000;
   assign mem[225055:225024] = 32'b11110110010010001001000111100000;
   assign mem[225087:225056] = 32'b11110110010110001011110111000000;
   assign mem[225119:225088] = 32'b00000001011100010011101010010000;
   assign mem[225151:225120] = 32'b11111100010111111001010101110100;
   assign mem[225183:225152] = 32'b00000100100100100111111101000000;
   assign mem[225215:225184] = 32'b11111110110011110001001100001110;
   assign mem[225247:225216] = 32'b00000011001100101011010111001100;
   assign mem[225279:225248] = 32'b00000010000110000000110111001000;
   assign mem[225311:225280] = 32'b11111111101010110101110101100100;
   assign mem[225343:225312] = 32'b11111010010111000000000101000000;
   assign mem[225375:225344] = 32'b11111011100110001110001001111000;
   assign mem[225407:225376] = 32'b00000000000100110001001000011001;
   assign mem[225439:225408] = 32'b00000101010110101001010011100000;
   assign mem[225471:225440] = 32'b00000011110000111000100101110100;
   assign mem[225503:225472] = 32'b11101101010100001011110110100000;
   assign mem[225535:225504] = 32'b11111011001011100001101110101000;
   assign mem[225567:225536] = 32'b00000100110110011111111100000000;
   assign mem[225599:225568] = 32'b00000101001111001000110110011000;
   assign mem[225631:225600] = 32'b11111001110111010111001111011000;
   assign mem[225663:225632] = 32'b11111001110001111011100001110000;
   assign mem[225695:225664] = 32'b11111100111111000000001100011000;
   assign mem[225727:225696] = 32'b00001110111100110000001011010000;
   assign mem[225759:225728] = 32'b11110000111100010100011001100000;
   assign mem[225791:225760] = 32'b00000111101111101110001111011000;
   assign mem[225823:225792] = 32'b11111011100100110000100010010000;
   assign mem[225855:225824] = 32'b11111000010111111010001000101000;
   assign mem[225887:225856] = 32'b11111001000100001101000110110000;
   assign mem[225919:225888] = 32'b00000101000010101101111110111000;
   assign mem[225951:225920] = 32'b00000000011111000110011001111011;
   assign mem[225983:225952] = 32'b11101000001010110100111100100000;
   assign mem[226015:225984] = 32'b11110101000101011100010000000000;
   assign mem[226047:226016] = 32'b11101110010100111110101000000000;
   assign mem[226079:226048] = 32'b00000110000011101011101111110000;
   assign mem[226111:226080] = 32'b11111111110001001001000110110011;
   assign mem[226143:226112] = 32'b11111100000011100010110000101100;
   assign mem[226175:226144] = 32'b11110110100100010010011010110000;
   assign mem[226207:226176] = 32'b00001011100001100001100111000000;
   assign mem[226239:226208] = 32'b00001000011111011001100011100000;
   assign mem[226271:226240] = 32'b11101000001111100110000110100000;
   assign mem[226303:226272] = 32'b11111101010101100110000011100000;
   assign mem[226335:226304] = 32'b11111111011011011100111101000101;
   assign mem[226367:226336] = 32'b00000000110101000011100011100010;
   assign mem[226399:226368] = 32'b11111111101000010111000110111001;
   assign mem[226431:226400] = 32'b00000011001111000010100000010000;
   assign mem[226463:226432] = 32'b11100010101001111110011100100000;
   assign mem[226495:226464] = 32'b00000010100010100010001010100000;
   assign mem[226527:226496] = 32'b11111100111100111011000011111000;
   assign mem[226559:226528] = 32'b00000010111001000101100110100100;
   assign mem[226591:226560] = 32'b11111000001110110111001010101000;
   assign mem[226623:226592] = 32'b00001001011000111011011111010000;
   assign mem[226655:226624] = 32'b00000100011100111100110110100000;
   assign mem[226687:226656] = 32'b00000001101000001010111110100100;
   assign mem[226719:226688] = 32'b11110111110110101010000000000000;
   assign mem[226751:226720] = 32'b00000010000101100000001011011000;
   assign mem[226783:226752] = 32'b11110111011010110111001010110000;
   assign mem[226815:226784] = 32'b00000111001100000010010000100000;
   assign mem[226847:226816] = 32'b11110010110111100001000101010000;
   assign mem[226879:226848] = 32'b11111001011100010000100110011000;
   assign mem[226911:226880] = 32'b00000000001010100011111110100011;
   assign mem[226943:226912] = 32'b11110010000010111010010110110000;
   assign mem[226975:226944] = 32'b11111010111100011001100010110000;
   assign mem[227007:226976] = 32'b11111010111000010011110111100000;
   assign mem[227039:227008] = 32'b00000100101010101101110101011000;
   assign mem[227071:227040] = 32'b00000010100011010001111001110100;
   assign mem[227103:227072] = 32'b11111110001011110111111011100010;
   assign mem[227135:227104] = 32'b11111010100111000100110001011000;
   assign mem[227167:227136] = 32'b00000010100100000000100101111100;
   assign mem[227199:227168] = 32'b00000000101100001111101100011100;
   assign mem[227231:227200] = 32'b11111110100001100011110111111000;
   assign mem[227263:227232] = 32'b00001001111101011000000010010000;
   assign mem[227295:227264] = 32'b00000011100010111100001011010000;
   assign mem[227327:227296] = 32'b00000111101111001111001000100000;
   assign mem[227359:227328] = 32'b11110111011011100111100110110000;
   assign mem[227391:227360] = 32'b11110011001111010111011000010000;
   assign mem[227423:227392] = 32'b00001011101101100011111011110000;
   assign mem[227455:227424] = 32'b00000000000110011101110110010010;
   assign mem[227487:227456] = 32'b11110101010110000001010100100000;
   assign mem[227519:227488] = 32'b11111011111111000001100100111000;
   assign mem[227551:227520] = 32'b00000000111000010100111010111010;
   assign mem[227583:227552] = 32'b00000100110111001110111011001000;
   assign mem[227615:227584] = 32'b11111000100111101101101101000000;
   assign mem[227647:227616] = 32'b00000111100010101001100001100000;
   assign mem[227679:227648] = 32'b11111100101100000001010111110000;
   assign mem[227711:227680] = 32'b11111010100001110001001011101000;
   assign mem[227743:227712] = 32'b00000010011010010101011100110100;
   assign mem[227775:227744] = 32'b00000100101011010001100001110000;
   assign mem[227807:227776] = 32'b11111001101001010001000000101000;
   assign mem[227839:227808] = 32'b11111010101101001110111001010000;
   assign mem[227871:227840] = 32'b11101001110101110101001000000000;
   assign mem[227903:227872] = 32'b11110110000000100101010011100000;
   assign mem[227935:227904] = 32'b00001000010010000100110001010000;
   assign mem[227967:227936] = 32'b00000010000100101001000011111100;
   assign mem[227999:227968] = 32'b11110001101111110100101010000000;
   assign mem[228031:228000] = 32'b11111111000001001100110101110010;
   assign mem[228063:228032] = 32'b11111001011011001101011011011000;
   assign mem[228095:228064] = 32'b00001101000110101110100101100000;
   assign mem[228127:228096] = 32'b11111100111111100101100010110000;
   assign mem[228159:228128] = 32'b00000001010111100001011111001000;
   assign mem[228191:228160] = 32'b00000011000110001010100001010100;
   assign mem[228223:228192] = 32'b00000000011001011010110010010011;
   assign mem[228255:228224] = 32'b11111011100000111110101110000000;
   assign mem[228287:228256] = 32'b11111010000100101011110110110000;
   assign mem[228319:228288] = 32'b11111101111011101110101110111000;
   assign mem[228351:228320] = 32'b00000010001011100101110001100000;
   assign mem[228383:228352] = 32'b00000011101000010100111011111000;
   assign mem[228415:228384] = 32'b11111110110100101000001111111110;
   assign mem[228447:228416] = 32'b11111001110101100110111101110000;
   assign mem[228479:228448] = 32'b11111111100101011110011010011011;
   assign mem[228511:228480] = 32'b00000000110111010010011010101111;
   assign mem[228543:228512] = 32'b00000000101010011011001000010011;
   assign mem[228575:228544] = 32'b00000111000000011111101101001000;
   assign mem[228607:228576] = 32'b11111111011001101101111010010110;
   assign mem[228639:228608] = 32'b11111101110110111100111010110000;
   assign mem[228671:228640] = 32'b11111001101011011100110101010000;
   assign mem[228703:228672] = 32'b11111000100101010000110110110000;
   assign mem[228735:228704] = 32'b00001000110001101101011010110000;
   assign mem[228767:228736] = 32'b11111101000100000110110110001000;
   assign mem[228799:228768] = 32'b11110111010101000111011100000000;
   assign mem[228831:228800] = 32'b11110101100011101000100001110000;
   assign mem[228863:228832] = 32'b11110110000000010010010000000000;
   assign mem[228895:228864] = 32'b11100101111110110110001011000000;
   assign mem[228927:228896] = 32'b11111100101111100000100110110000;
   assign mem[228959:228928] = 32'b00000110011110011111000100110000;
   assign mem[228991:228960] = 32'b11111111111000010101111101000100;
   assign mem[229023:228992] = 32'b11110111101101000000100001010000;
   assign mem[229055:229024] = 32'b11111110100000011110111101101100;
   assign mem[229087:229056] = 32'b00000101101110100001001100010000;
   assign mem[229119:229088] = 32'b00001001011101010110000000010000;
   assign mem[229151:229120] = 32'b11110110111111100111011001100000;
   assign mem[229183:229152] = 32'b11110000100101011111111011010000;
   assign mem[229215:229184] = 32'b00000100010011110110100100011000;
   assign mem[229247:229216] = 32'b11111000011010011101011000001000;
   assign mem[229279:229248] = 32'b00000100010110010110100001000000;
   assign mem[229311:229280] = 32'b11111111111100111000001110000110;
   assign mem[229343:229312] = 32'b11111000110111101101111111110000;
   assign mem[229375:229344] = 32'b11111001101101000110010111111000;
   assign mem[229407:229376] = 32'b00000100011010001101110110010000;
   assign mem[229439:229408] = 32'b00000100110111101000110000111000;
   assign mem[229471:229440] = 32'b11111001000000011011001111000000;
   assign mem[229503:229472] = 32'b11111011010101000111010010101000;
   assign mem[229535:229504] = 32'b00000000000111011100110001010011;
   assign mem[229567:229536] = 32'b11111011100001001101000101110000;
   assign mem[229599:229568] = 32'b00000000100111110010010010011011;
   assign mem[229631:229600] = 32'b11111011001011111100010000100000;
   assign mem[229663:229632] = 32'b00000010101000101111001001010100;
   assign mem[229695:229664] = 32'b11111110111001101010101011000110;
   assign mem[229727:229696] = 32'b00001010001011100100101011110000;
   assign mem[229759:229728] = 32'b11111101101010100101101110111100;
   assign mem[229791:229760] = 32'b00000010100100000101100000110000;
   assign mem[229823:229792] = 32'b11111000101001111100100010100000;
   assign mem[229855:229824] = 32'b11111100001110110101000101001000;
   assign mem[229887:229856] = 32'b11101111101011001010000010100000;
   assign mem[229919:229888] = 32'b00000100110001100101111000100000;
   assign mem[229951:229920] = 32'b00000110110001001001110010101000;
   assign mem[229983:229952] = 32'b00000000001001100010111100111011;
   assign mem[230015:229984] = 32'b11101111111000101000011101100000;
   assign mem[230047:230016] = 32'b00001000101001110111110000000000;
   assign mem[230079:230048] = 32'b00000111000001011001010101110000;
   assign mem[230111:230080] = 32'b00000101011001111010001110110000;
   assign mem[230143:230112] = 32'b00000001100011111001000101101110;
   assign mem[230175:230144] = 32'b11111110001111110111111101111100;
   assign mem[230207:230176] = 32'b11111111001010000101010110111111;
   assign mem[230239:230208] = 32'b00000010111011111000110000100100;
   assign mem[230271:230240] = 32'b00000010001001011000010011101100;
   assign mem[230303:230272] = 32'b11111110011011100100101011011010;
   assign mem[230335:230304] = 32'b11111111001010011101000100000000;
   assign mem[230367:230336] = 32'b00000011100000001011111101010000;
   assign mem[230399:230368] = 32'b11111110010000001000111100010000;
   assign mem[230431:230400] = 32'b11110110010001100101001000000000;
   assign mem[230463:230432] = 32'b00000001001101001110011001001100;
   assign mem[230495:230464] = 32'b00000000101110000111110101000010;
   assign mem[230527:230496] = 32'b11111111101110001111010011010100;
   assign mem[230559:230528] = 32'b11111111111100110100100100111001;
   assign mem[230591:230560] = 32'b00000011010000000111101110000000;
   assign mem[230623:230592] = 32'b11110101100100000001000111010000;
   assign mem[230655:230624] = 32'b00000111111100000110110000011000;
   assign mem[230687:230656] = 32'b11110111000001011100110001000000;
   assign mem[230719:230688] = 32'b11111111001000011011111110001111;
   assign mem[230751:230720] = 32'b11111100100111001111111101111000;
   assign mem[230783:230752] = 32'b11111001111011001011100110100000;
   assign mem[230815:230784] = 32'b11111000100100101100110101010000;
   assign mem[230847:230816] = 32'b11111000000110011111100000010000;
   assign mem[230879:230848] = 32'b00000100101100000011011001100000;
   assign mem[230911:230880] = 32'b00000000110101000010010110100011;
   assign mem[230943:230912] = 32'b00000101011000010011010010111000;
   assign mem[230975:230944] = 32'b00000000111010001100010110110100;
   assign mem[231007:230976] = 32'b00000011110111011011101000011100;
   assign mem[231039:231008] = 32'b00000011101100101110111110111000;
   assign mem[231071:231040] = 32'b00000000010011100010011111101101;
   assign mem[231103:231072] = 32'b00000010111111101011110111101000;
   assign mem[231135:231104] = 32'b11111101000010100110100011111100;
   assign mem[231167:231136] = 32'b11111101100010010010111110010000;
   assign mem[231199:231168] = 32'b00000101110101100111101010100000;
   assign mem[231231:231200] = 32'b00000010110110111010011010000100;
   assign mem[231263:231232] = 32'b00000000101010000100110101001101;
   assign mem[231295:231264] = 32'b11111111001001001010010010111011;
   assign mem[231327:231296] = 32'b11110100011001001000010100010000;
   assign mem[231359:231328] = 32'b00000100110100101100001010100000;
   assign mem[231391:231360] = 32'b00000001101001011011001111001000;
   assign mem[231423:231392] = 32'b00000010001101111011010111010100;
   assign mem[231455:231424] = 32'b00000111111101000000110000000000;
   assign mem[231487:231456] = 32'b11111100010001000001111100011100;
   assign mem[231519:231488] = 32'b11111010101010011001001011110000;
   assign mem[231551:231520] = 32'b11111000011101000011001000111000;
   assign mem[231583:231552] = 32'b11111011001111100011001001111000;
   assign mem[231615:231584] = 32'b00000001000000101000111100010000;
   assign mem[231647:231616] = 32'b00000101110011001111011000000000;
   assign mem[231679:231648] = 32'b11111000111000010101110011101000;
   assign mem[231711:231680] = 32'b00000010010010011000101001000100;
   assign mem[231743:231712] = 32'b11111111011110101011011010101010;
   assign mem[231775:231744] = 32'b11111010011110101010011110000000;
   assign mem[231807:231776] = 32'b11110100011101110101111011110000;
   assign mem[231839:231808] = 32'b00000011010010110001000101111000;
   assign mem[231871:231840] = 32'b00000001111011101111001101000000;
   assign mem[231903:231872] = 32'b00000010010000101001100101111100;
   assign mem[231935:231904] = 32'b00000100001010000011111000110000;
   assign mem[231967:231936] = 32'b00000010011010101010100100010000;
   assign mem[231999:231968] = 32'b00000010100111000101100111101100;
   assign mem[232031:232000] = 32'b11111011101010100010110100101000;
   assign mem[232063:232032] = 32'b11111010001011110010000011011000;
   assign mem[232095:232064] = 32'b00001001011011100000101000010000;
   assign mem[232127:232096] = 32'b11111101000100001000101110111100;
   assign mem[232159:232128] = 32'b11111001101000111111110111010000;
   assign mem[232191:232160] = 32'b11111001010110010010100000011000;
   assign mem[232223:232192] = 32'b11111011110110001111001101110000;
   assign mem[232255:232224] = 32'b00000110001011111011111110010000;
   assign mem[232287:232256] = 32'b00000010000100101010001010010000;
   assign mem[232319:232288] = 32'b11111100111001101101001001100000;
   assign mem[232351:232320] = 32'b11111110110000001101001011100110;
   assign mem[232383:232352] = 32'b00000001101000011011010001110010;
   assign mem[232415:232384] = 32'b11110111001011111001101111000000;
   assign mem[232447:232416] = 32'b11111101010101111001001011010100;
   assign mem[232479:232448] = 32'b00001010001010101100011100000000;
   assign mem[232511:232480] = 32'b11110101010101011001000011010000;
   assign mem[232543:232512] = 32'b11111101110011000110101100001100;
   assign mem[232575:232544] = 32'b11111111000111111000111011110111;
   assign mem[232607:232576] = 32'b00000011001100000100011101011000;
   assign mem[232639:232608] = 32'b00000001000000111110010100001100;
   assign mem[232671:232640] = 32'b00000001011001100111000110110100;
   assign mem[232703:232672] = 32'b11101001000011110011110100100000;
   assign mem[232735:232704] = 32'b11101000011001010110100011000000;
   assign mem[232767:232736] = 32'b11111000011011000011001001100000;
   assign mem[232799:232768] = 32'b00000011111111011100011100100000;
   assign mem[232831:232800] = 32'b00000011100010101010000011110000;
   assign mem[232863:232832] = 32'b00000001100110011110111111100110;
   assign mem[232895:232864] = 32'b11111010100010001011001011010000;
   assign mem[232927:232896] = 32'b00000101101000111110011111101000;
   assign mem[232959:232928] = 32'b00001001000111111000101100100000;
   assign mem[232991:232960] = 32'b00000010000111110010111100000100;
   assign mem[233023:232992] = 32'b11100101010100000100010110100000;
   assign mem[233055:233024] = 32'b11101111110101111101110001100000;
   assign mem[233087:233056] = 32'b11111010100100111011010011110000;
   assign mem[233119:233088] = 32'b00000110011001101111000101110000;
   assign mem[233151:233120] = 32'b00000100001011111101001100000000;
   assign mem[233183:233152] = 32'b00000001000101111011100011110100;
   assign mem[233215:233184] = 32'b00000001100011110001101011110110;
   assign mem[233247:233216] = 32'b00001000100111011110000111110000;
   assign mem[233279:233248] = 32'b00000101000110111010001001000000;
   assign mem[233311:233280] = 32'b11111111111011001000100101011100;
   assign mem[233343:233312] = 32'b00000001101100101110001010110010;
   assign mem[233375:233344] = 32'b11110110011101101011001110000000;
   assign mem[233407:233376] = 32'b11111001100110101111001011000000;
   assign mem[233439:233408] = 32'b00000101000010110000100001100000;
   assign mem[233471:233440] = 32'b11110001000110000101011000010000;
   assign mem[233503:233472] = 32'b00000110110001011000100110100000;
   assign mem[233535:233504] = 32'b00001101111001010011101110000000;
   assign mem[233567:233536] = 32'b11111011001100111100100110110000;
   assign mem[233599:233568] = 32'b00000000110010000101111100011010;
   assign mem[233631:233600] = 32'b00000011011111010110101101000000;
   assign mem[233663:233632] = 32'b11111011000100111010100101100000;
   assign mem[233695:233664] = 32'b11101010100001010100000110000000;
   assign mem[233727:233696] = 32'b11111010001111101011000101010000;
   assign mem[233759:233728] = 32'b00000001011111001110010011100110;
   assign mem[233791:233760] = 32'b00000100001101000000101010100000;
   assign mem[233823:233792] = 32'b00000000111010101101010100010111;
   assign mem[233855:233824] = 32'b11111111011000010100001001101011;
   assign mem[233887:233856] = 32'b00001001010101100000011101010000;
   assign mem[233919:233888] = 32'b00000000111110011101010100000101;
   assign mem[233951:233920] = 32'b00000011111100111000000001010000;
   assign mem[233983:233952] = 32'b00000110100100100010011100110000;
   assign mem[234015:233984] = 32'b00000100001011110010101000101000;
   assign mem[234047:234016] = 32'b11111111000100111010111110001110;
   assign mem[234079:234048] = 32'b00000011001011010111100111010000;
   assign mem[234111:234080] = 32'b11111011110110000010000000000000;
   assign mem[234143:234112] = 32'b00000111110000101001100000010000;
   assign mem[234175:234144] = 32'b00000111000000101100011101110000;
   assign mem[234207:234176] = 32'b11111101100000111101111100000000;
   assign mem[234239:234208] = 32'b11111010100101010010000011010000;
   assign mem[234271:234240] = 32'b11111100110111111100111011110000;
   assign mem[234303:234272] = 32'b11111110111111101110111000100110;
   assign mem[234335:234304] = 32'b00001001100110100000011010010000;
   assign mem[234367:234336] = 32'b11110011001110000000010100110000;
   assign mem[234399:234368] = 32'b00000000101110001111100000011101;
   assign mem[234431:234400] = 32'b00000110000011100011100001001000;
   assign mem[234463:234432] = 32'b11111110100110100001100000000000;
   assign mem[234495:234464] = 32'b11110101001011101111101010000000;
   assign mem[234527:234496] = 32'b00000101101110010101111001010000;
   assign mem[234559:234528] = 32'b00000111000001001010100100011000;
   assign mem[234591:234560] = 32'b11110001111111101111101000010000;
   assign mem[234623:234592] = 32'b11110100010110010111011100110000;
   assign mem[234655:234624] = 32'b00001001110000110101011000000000;
   assign mem[234687:234656] = 32'b00000100010110100110100101001000;
   assign mem[234719:234688] = 32'b11111001101101110010010110001000;
   assign mem[234751:234720] = 32'b11110111100001011011011010100000;
   assign mem[234783:234752] = 32'b11111111111011000001000110011111;
   assign mem[234815:234784] = 32'b00001111101111110101001111100000;
   assign mem[234847:234816] = 32'b11111011100100010110100101110000;
   assign mem[234879:234848] = 32'b11110111000001101001101011010000;
   assign mem[234911:234880] = 32'b00000011110010100010010000010100;
   assign mem[234943:234912] = 32'b11101100101111111100011011100000;
   assign mem[234975:234944] = 32'b11110011011111101100110011010000;
   assign mem[235007:234976] = 32'b11111100101111011001011001111000;
   assign mem[235039:235008] = 32'b11111111101101111001110110110100;
   assign mem[235071:235040] = 32'b11111111100001000111110001000011;
   assign mem[235103:235072] = 32'b00000100011101100110010001011000;
   assign mem[235135:235104] = 32'b00001010101001001111101110010000;
   assign mem[235167:235136] = 32'b00000000110001010110011000001010;
   assign mem[235199:235168] = 32'b00000010010110000011101111011100;
   assign mem[235231:235200] = 32'b11110010011010000001111000000000;
   assign mem[235263:235232] = 32'b11111100110101000000010101001000;
   assign mem[235295:235264] = 32'b11111101101111101101000001111100;
   assign mem[235327:235296] = 32'b11111101101100111010100010010000;
   assign mem[235359:235328] = 32'b00000110001011110010110001110000;
   assign mem[235391:235360] = 32'b00000001111010111010101000110000;
   assign mem[235423:235392] = 32'b11100100110110000110101001000000;
   assign mem[235455:235424] = 32'b00000110101000001000110110011000;
   assign mem[235487:235456] = 32'b11111100010011110010011000110100;
   assign mem[235519:235488] = 32'b00000101010110100110001000100000;
   assign mem[235551:235520] = 32'b00000000110010111100010101011100;
   assign mem[235583:235552] = 32'b00000001101000111111100110101000;
   assign mem[235615:235584] = 32'b11111010010111111100100011011000;
   assign mem[235647:235616] = 32'b11111111000101101111100000010111;
   assign mem[235679:235648] = 32'b00000010100111010001100000001000;
   assign mem[235711:235680] = 32'b11111010111101101101111010101000;
   assign mem[235743:235712] = 32'b00000000011010010111011101010111;
   assign mem[235775:235744] = 32'b00000010111001011110101000101100;
   assign mem[235807:235776] = 32'b11111100011010100011010111111100;
   assign mem[235839:235808] = 32'b11111101011111100110010011000000;
   assign mem[235871:235840] = 32'b00000100101111100100110010000000;
   assign mem[235903:235872] = 32'b11111101110010011000001100110100;
   assign mem[235935:235904] = 32'b11111100110101011101101100011000;
   assign mem[235967:235936] = 32'b11111000010010010100100111110000;
   assign mem[235999:235968] = 32'b00000011000110000101011001011000;
   assign mem[236031:236000] = 32'b11111110100001100000000000111010;
   assign mem[236063:236032] = 32'b00000010111000000000111000010100;
   assign mem[236095:236064] = 32'b11111101101000010010001101001100;
   assign mem[236127:236096] = 32'b11111101110111011011000101111000;
   assign mem[236159:236128] = 32'b00000110111111000101000100000000;
   assign mem[236191:236160] = 32'b11111010010111010101011111001000;
   assign mem[236223:236192] = 32'b11110000100000101010111001000000;
   assign mem[236255:236224] = 32'b00000001010011101000011011110100;
   assign mem[236287:236256] = 32'b11110100111100011000010011000000;
   assign mem[236319:236288] = 32'b00000111011010001111100001000000;
   assign mem[236351:236320] = 32'b00000001101011101100101011011010;
   assign mem[236383:236352] = 32'b11110111000111001000110001010000;
   assign mem[236415:236384] = 32'b00000001100101000000110101111100;
   assign mem[236447:236416] = 32'b00000101000010001011001000100000;
   assign mem[236479:236448] = 32'b00001000011100101100010111110000;
   assign mem[236511:236480] = 32'b11111001100001110011110110010000;
   assign mem[236543:236512] = 32'b00000010000110011110011010101100;
   assign mem[236575:236544] = 32'b00000100011101110111000111100000;
   assign mem[236607:236576] = 32'b00001000011110110000000111000000;
   assign mem[236639:236608] = 32'b11111100000011010011000111101000;
   assign mem[236671:236640] = 32'b11101111010110000100111011100000;
   assign mem[236703:236672] = 32'b00001011001000111011100111010000;
   assign mem[236735:236704] = 32'b11111110111010010100011010111110;
   assign mem[236767:236736] = 32'b11110010111001001111010100110000;
   assign mem[236799:236768] = 32'b11111011110100000100100011001000;
   assign mem[236831:236800] = 32'b11110110111000100000001110100000;
   assign mem[236863:236832] = 32'b11111001001000001000000111011000;
   assign mem[236895:236864] = 32'b00000010100101001010101111000000;
   assign mem[236927:236896] = 32'b11111101101000011001101110101100;
   assign mem[236959:236928] = 32'b00000011011110000101011001101100;
   assign mem[236991:236960] = 32'b11111110011100111001001011000110;
   assign mem[237023:236992] = 32'b11111011010010101111100000100000;
   assign mem[237055:237024] = 32'b00000011100001110010100111011000;
   assign mem[237087:237056] = 32'b11111100010010110001100000011000;
   assign mem[237119:237088] = 32'b00000010100111100110111100001100;
   assign mem[237151:237120] = 32'b00000011101010011100000111011100;
   assign mem[237183:237152] = 32'b11111101010111010010101000010100;
   assign mem[237215:237184] = 32'b00000001000001000011010100011010;
   assign mem[237247:237216] = 32'b00000001010001111111010011101100;
   assign mem[237279:237248] = 32'b11111101111010000101101011000000;
   assign mem[237311:237280] = 32'b00000011100101111100110011010100;
   assign mem[237343:237312] = 32'b11111110001001011011111111000110;
   assign mem[237375:237344] = 32'b00000011000111101101110101000000;
   assign mem[237407:237376] = 32'b11111100101011101110011101000000;
   assign mem[237439:237408] = 32'b00000001110101111100010111011010;
   assign mem[237471:237440] = 32'b00000011011111001000101000011100;
   assign mem[237503:237472] = 32'b11101111111000111011110110100000;
   assign mem[237535:237504] = 32'b11111001010001001011001110000000;
   assign mem[237567:237536] = 32'b11110110111111101000000000000000;
   assign mem[237599:237568] = 32'b00000110011011011011111001110000;
   assign mem[237631:237600] = 32'b00001000101111101111110010000000;
   assign mem[237663:237632] = 32'b00000110100110011011111001101000;
   assign mem[237695:237664] = 32'b11111001000110001110101001011000;
   assign mem[237727:237696] = 32'b00000011001010111110011111101100;
   assign mem[237759:237728] = 32'b00001000010110010101111000110000;
   assign mem[237791:237760] = 32'b11110101100010000000101100000000;
   assign mem[237823:237792] = 32'b00000100010101011101110101010000;
   assign mem[237855:237824] = 32'b00001001000000110001111100010000;
   assign mem[237887:237856] = 32'b00000010001101100010000101100100;
   assign mem[237919:237888] = 32'b11101111111001000110011101000000;
   assign mem[237951:237920] = 32'b11111100100110101111110001010100;
   assign mem[237983:237952] = 32'b11110010110100011100001010110000;
   assign mem[238015:237984] = 32'b00001010011001010011101001000000;
   assign mem[238047:238016] = 32'b11111010100101100101110100001000;
   assign mem[238079:238048] = 32'b11110001101100000111001000010000;
   assign mem[238111:238080] = 32'b00000000110111000110011001101110;
   assign mem[238143:238112] = 32'b00000000100010110010100110101110;
   assign mem[238175:238144] = 32'b11110011101100010000000011000000;
   assign mem[238207:238176] = 32'b11110001100101110010010001000000;
   assign mem[238239:238208] = 32'b00000100100100110001111110110000;
   assign mem[238271:238240] = 32'b00000100110000010010100111000000;
   assign mem[238303:238272] = 32'b11110110111110110000000010000000;
   assign mem[238335:238304] = 32'b00000010011000111101000000110000;
   assign mem[238367:238336] = 32'b00000111110010111101010001101000;
   assign mem[238399:238368] = 32'b00001010000101011100011000110000;
   assign mem[238431:238400] = 32'b11111010001000110101100100111000;
   assign mem[238463:238432] = 32'b00000011011110000001101100001000;
   assign mem[238495:238464] = 32'b00000101001111100101100000001000;
   assign mem[238527:238496] = 32'b00000011101010011111001001010100;
   assign mem[238559:238528] = 32'b11111001000111111111011110010000;
   assign mem[238591:238560] = 32'b00000110101101101001100111111000;
   assign mem[238623:238592] = 32'b11111000101111001100010111000000;
   assign mem[238655:238624] = 32'b00001000000110111010010100000000;
   assign mem[238687:238656] = 32'b11110001110011000111100011100000;
   assign mem[238719:238688] = 32'b11110111011001001001000010110000;
   assign mem[238751:238720] = 32'b11100101001110111101010001000000;
   assign mem[238783:238752] = 32'b00000011000010010010000011000100;
   assign mem[238815:238784] = 32'b00000011010001001011110001111100;
   assign mem[238847:238816] = 32'b00000101110000110010101100001000;
   assign mem[238879:238848] = 32'b00000101000011101010000100000000;
   assign mem[238911:238880] = 32'b00000100110011001101000111001000;
   assign mem[238943:238912] = 32'b11011011010101111100101111000000;
   assign mem[238975:238944] = 32'b00000011100001110110010001100100;
   assign mem[239007:238976] = 32'b11111010010000110101110000101000;
   assign mem[239039:239008] = 32'b00000010001101101100101101101000;
   assign mem[239071:239040] = 32'b00000010101011100101000111110000;
   assign mem[239103:239072] = 32'b11111101101010001110101100001000;
   assign mem[239135:239104] = 32'b11110001000000100100101010100000;
   assign mem[239167:239136] = 32'b11111110100000010100010100011110;
   assign mem[239199:239168] = 32'b00000101001000000111001101010000;
   assign mem[239231:239200] = 32'b00000000110111011100111101001101;
   assign mem[239263:239232] = 32'b00000110000011010101001100000000;
   assign mem[239295:239264] = 32'b11111111001101101000001000100011;
   assign mem[239327:239296] = 32'b11111101000011110101110111010100;
   assign mem[239359:239328] = 32'b00000001101000011111111010111110;
   assign mem[239391:239360] = 32'b00000010110100001010001001101100;
   assign mem[239423:239392] = 32'b11101101111100010110001010000000;
   assign mem[239455:239424] = 32'b11111101111000100101011011010100;
   assign mem[239487:239456] = 32'b11110111010010000110100000110000;
   assign mem[239519:239488] = 32'b00000101101101010011010100011000;
   assign mem[239551:239520] = 32'b00000010110101100010100001101000;
   assign mem[239583:239552] = 32'b00000100101001100000110011000000;
   assign mem[239615:239584] = 32'b11110001001110101111001011010000;
   assign mem[239647:239616] = 32'b00000111101011001110110011110000;
   assign mem[239679:239648] = 32'b00000110110111010100111110010000;
   assign mem[239711:239680] = 32'b00000011100011001100011101010000;
   assign mem[239743:239712] = 32'b11111100000000000101001110011000;
   assign mem[239775:239744] = 32'b11111010010100000110111010011000;
   assign mem[239807:239776] = 32'b11111101100100001110100110011100;
   assign mem[239839:239808] = 32'b11111111001000011100000111111110;
   assign mem[239871:239840] = 32'b11111011010000010101100110010000;
   assign mem[239903:239872] = 32'b00000011010010010110001011000000;
   assign mem[239935:239904] = 32'b00000100011110111111111111111000;
   assign mem[239967:239936] = 32'b00000011011101011100101101001100;
   assign mem[239999:239968] = 32'b00000000011001111111110000010011;
   assign mem[240031:240000] = 32'b00000011010101000110111000010100;
   assign mem[240063:240032] = 32'b00000001000001011001101000011100;
   assign mem[240095:240064] = 32'b11110111111100111101010110110000;
   assign mem[240127:240096] = 32'b11110111010100011110100001010000;
   assign mem[240159:240128] = 32'b11111110010011011001011111010100;
   assign mem[240191:240160] = 32'b00000000100000111000101111000111;
   assign mem[240223:240192] = 32'b00000000111111010100111111110000;
   assign mem[240255:240224] = 32'b11111010110100101010010011100000;
   assign mem[240287:240256] = 32'b00000100111011011001001011101000;
   assign mem[240319:240288] = 32'b00000100110111101001010111010000;
   assign mem[240351:240320] = 32'b00000001001110101110000111110110;
   assign mem[240383:240352] = 32'b11111101110011001100101011010000;
   assign mem[240415:240384] = 32'b11111111010110111001110010011100;
   assign mem[240447:240416] = 32'b11111101011111111110010111111000;
   assign mem[240479:240448] = 32'b11111100010001011001110111001000;
   assign mem[240511:240480] = 32'b00000011101000011110001011101100;
   assign mem[240543:240512] = 32'b11111100110010010000000010011000;
   assign mem[240575:240544] = 32'b11111110100101110001100110101000;
   assign mem[240607:240576] = 32'b11111101010101101110011101011100;
   assign mem[240639:240608] = 32'b11111100010000000101111000110000;
   assign mem[240671:240640] = 32'b00000011101110101010010110101000;
   assign mem[240703:240672] = 32'b11111101001010100100100001000100;
   assign mem[240735:240704] = 32'b00000110000100110010111000101000;
   assign mem[240767:240736] = 32'b11101100011001101100110101000000;
   assign mem[240799:240768] = 32'b00000100000000001011010000000000;
   assign mem[240831:240800] = 32'b00000100101001011100111110110000;
   assign mem[240863:240832] = 32'b00000000000010110001000110110010;
   assign mem[240895:240864] = 32'b00000100000010100100010110100000;
   assign mem[240927:240896] = 32'b11111100000111000101100001001000;
   assign mem[240959:240928] = 32'b11111111110101101101001100110101;
   assign mem[240991:240960] = 32'b00000100010010011001100101001000;
   assign mem[241023:240992] = 32'b00000001101101101011101000100010;
   assign mem[241055:241024] = 32'b00000011001001101101011101110000;
   assign mem[241087:241056] = 32'b11111011001111010010110100100000;
   assign mem[241119:241088] = 32'b00000101010010011111000001101000;
   assign mem[241151:241120] = 32'b11111110011110101011111001111110;
   assign mem[241183:241152] = 32'b00000100100101011010010000000000;
   assign mem[241215:241184] = 32'b11111101101000001011011001110000;
   assign mem[241247:241216] = 32'b00000000100111110101100000001110;
   assign mem[241279:241248] = 32'b11111101001011010010101100101000;
   assign mem[241311:241280] = 32'b00000101100110100001000001110000;
   assign mem[241343:241312] = 32'b00000001000001101010100000110000;
   assign mem[241375:241344] = 32'b00000010000101101011100011010000;
   assign mem[241407:241376] = 32'b11110101011111001111111010100000;
   assign mem[241439:241408] = 32'b00000001010110100110010010010100;
   assign mem[241471:241440] = 32'b00000000111100010010011101011101;
   assign mem[241503:241472] = 32'b11111010100010001110111000001000;
   assign mem[241535:241504] = 32'b11111101110011000011000110001100;
   assign mem[241567:241536] = 32'b00001000010111010001000110110000;
   assign mem[241599:241568] = 32'b11111101000101010001001111001100;
   assign mem[241631:241600] = 32'b11111011111000011000001010100000;
   assign mem[241663:241632] = 32'b11111111011000101100100111001000;
   assign mem[241695:241664] = 32'b00000000110011100010101100110111;
   assign mem[241727:241696] = 32'b00000101000001000110110000010000;
   assign mem[241759:241728] = 32'b11111110101101111011111010010000;
   assign mem[241791:241760] = 32'b00000001110101100001010010100110;
   assign mem[241823:241792] = 32'b11111100111001101110101011010100;
   assign mem[241855:241824] = 32'b11111101101101001100010100000000;
   assign mem[241887:241856] = 32'b00000001000000001111000000001000;
   assign mem[241919:241888] = 32'b00000000111001111110000010001111;
   assign mem[241951:241920] = 32'b11110110111101100011010110000000;
   assign mem[241983:241952] = 32'b11110111000101001011000101010000;
   assign mem[242015:241984] = 32'b00000010100111110000001010100100;
   assign mem[242047:242016] = 32'b11111111110101100110100011110110;
   assign mem[242079:242048] = 32'b00000100111010100101100111000000;
   assign mem[242111:242080] = 32'b00000000101001110011010111111011;
   assign mem[242143:242112] = 32'b11110110101000011001111000010000;
   assign mem[242175:242144] = 32'b00000010110111000101101111101000;
   assign mem[242207:242176] = 32'b11111011010001110010111011111000;
   assign mem[242239:242208] = 32'b00000010100000110010101001101000;
   assign mem[242271:242240] = 32'b11111010101100011100100101110000;
   assign mem[242303:242272] = 32'b11110101000010101001101001010000;
   assign mem[242335:242304] = 32'b00000011111001101001110001101100;
   assign mem[242367:242336] = 32'b11110101101101001100010001000000;
   assign mem[242399:242368] = 32'b00000100110110000011101010100000;
   assign mem[242431:242400] = 32'b11111011101011001011011100111000;
   assign mem[242463:242432] = 32'b11101100000011111000001111100000;
   assign mem[242495:242464] = 32'b11111100000111010011001110000100;
   assign mem[242527:242496] = 32'b00000010100001011101010011011100;
   assign mem[242559:242528] = 32'b00000100011100001001101101010000;
   assign mem[242591:242560] = 32'b11111010100111101011100011011000;
   assign mem[242623:242592] = 32'b11111101000010001011100101011000;
   assign mem[242655:242624] = 32'b11111010111110111101001110011000;
   assign mem[242687:242656] = 32'b11111111001100001100100000010111;
   assign mem[242719:242688] = 32'b00000110011011101011100000000000;
   assign mem[242751:242720] = 32'b00000011100111111001001101100100;
   assign mem[242783:242752] = 32'b11110101000001011011110101100000;
   assign mem[242815:242784] = 32'b00000101110101110001100100000000;
   assign mem[242847:242816] = 32'b11111000001011011000010011110000;
   assign mem[242879:242848] = 32'b00000000100111000000000101000101;
   assign mem[242911:242880] = 32'b11111100100101011000101010001100;
   assign mem[242943:242912] = 32'b00000000010111000011000011110100;
   assign mem[242975:242944] = 32'b11110010011111010010010010110000;
   assign mem[243007:242976] = 32'b00010001000000010100000111100000;
   assign mem[243039:243008] = 32'b11111100100110000000101001110100;
   assign mem[243071:243040] = 32'b11111011011101010001111001000000;
   assign mem[243103:243072] = 32'b00000011010001011001100010011100;
   assign mem[243135:243104] = 32'b11111100111000011001101100111100;
   assign mem[243167:243136] = 32'b11111011001101001000110010001000;
   assign mem[243199:243168] = 32'b00000111010011110101111100101000;
   assign mem[243231:243200] = 32'b00000100001101100000110000000000;
   assign mem[243263:243232] = 32'b11111101110101011110100000011100;
   assign mem[243295:243264] = 32'b11110101001101100111101111010000;
   assign mem[243327:243296] = 32'b11111010111010100010010100101000;
   assign mem[243359:243328] = 32'b00001000110111001111001111010000;
   assign mem[243391:243360] = 32'b11111011110011100011110000000000;
   assign mem[243423:243392] = 32'b00000001000010000110101100101010;
   assign mem[243455:243424] = 32'b00001011000101011100100111000000;
   assign mem[243487:243456] = 32'b11111011011000100100010010000000;
   assign mem[243519:243488] = 32'b11111001100101100101111000001000;
   assign mem[243551:243520] = 32'b11101010010110110011010010100000;
   assign mem[243583:243552] = 32'b11111110111100011110111100101010;
   assign mem[243615:243584] = 32'b11111000001101000101100000101000;
   assign mem[243647:243616] = 32'b11111101011010010100010011110100;
   assign mem[243679:243648] = 32'b00000101100100001001110110000000;
   assign mem[243711:243680] = 32'b00000000011101000011001010100001;
   assign mem[243743:243712] = 32'b11101000101110000010011010000000;
   assign mem[243775:243744] = 32'b00000010010010001111111011001100;
   assign mem[243807:243776] = 32'b00000101011100001101001011101000;
   assign mem[243839:243808] = 32'b00000111110100000101100111100000;
   assign mem[243871:243840] = 32'b11111000000010011101000010001000;
   assign mem[243903:243872] = 32'b11110111001101100010011101100000;
   assign mem[243935:243904] = 32'b00000100101101101001000001100000;
   assign mem[243967:243936] = 32'b11111110010000000101001011011110;
   assign mem[243999:243968] = 32'b11111101110011110010011011011000;
   assign mem[244031:244000] = 32'b11111101011010011001011101110100;
   assign mem[244063:244032] = 32'b11111110011110111101101101010110;
   assign mem[244095:244064] = 32'b00000011010110000001111011100000;
   assign mem[244127:244096] = 32'b00000000001111110000011000010111;
   assign mem[244159:244128] = 32'b11111100001101101000000000000000;
   assign mem[244191:244160] = 32'b00000000010111110000010011000101;
   assign mem[244223:244192] = 32'b11111001000011110100000110100000;
   assign mem[244255:244224] = 32'b00000001100011101001010101010010;
   assign mem[244287:244256] = 32'b11110111100011110011000010000000;
   assign mem[244319:244288] = 32'b00000011101101110111110110010000;
   assign mem[244351:244320] = 32'b11111111011011011011100111000111;
   assign mem[244383:244352] = 32'b00000110001111010000001010010000;
   assign mem[244415:244384] = 32'b00000100001000100010000001110000;
   assign mem[244447:244416] = 32'b11111111101101001101000110010010;
   assign mem[244479:244448] = 32'b11111111101110000010011111101010;
   assign mem[244511:244480] = 32'b00000001110100001010011100000010;
   assign mem[244543:244512] = 32'b00000101111110011101101100001000;
   assign mem[244575:244544] = 32'b00000101010001000011101000100000;
   assign mem[244607:244576] = 32'b00000100001100111011010111101000;
   assign mem[244639:244608] = 32'b11111110110110010111011010000000;
   assign mem[244671:244640] = 32'b11111011111111011000010000001000;
   assign mem[244703:244672] = 32'b11111101101110110000001000110000;
   assign mem[244735:244704] = 32'b00001100000101010011111010000000;
   assign mem[244767:244736] = 32'b11111110111110000101010101101110;
   assign mem[244799:244768] = 32'b11101101001001010110111110000000;
   assign mem[244831:244800] = 32'b00000100001011100000100111000000;
   assign mem[244863:244832] = 32'b11111101111001000110001100110000;
   assign mem[244895:244864] = 32'b00000000111111011010010110000010;
   assign mem[244927:244896] = 32'b11110100000010000001001111110000;
   assign mem[244959:244928] = 32'b00000100100011111001110101110000;
   assign mem[244991:244960] = 32'b11111110011011000000010000000110;
   assign mem[245023:244992] = 32'b00000001111000011010110111010110;
   assign mem[245055:245024] = 32'b11111101011101100001011010101100;
   assign mem[245087:245056] = 32'b11111011011010010100000100000000;
   assign mem[245119:245088] = 32'b00000011001000100010111000001000;
   assign mem[245151:245120] = 32'b00000000011100110110001110110100;
   assign mem[245183:245152] = 32'b00000001000010101001100101000000;
   assign mem[245215:245184] = 32'b11111100001000011100010110100000;
   assign mem[245247:245216] = 32'b11111011000000110110100101111000;
   assign mem[245279:245248] = 32'b11111110111000010111001001001000;
   assign mem[245311:245280] = 32'b00000011011110011110101001101000;
   assign mem[245343:245312] = 32'b00000110011000010011000011110000;
   assign mem[245375:245344] = 32'b00000000101100101100001010001111;
   assign mem[245407:245376] = 32'b11111110101011100001110100111110;
   assign mem[245439:245408] = 32'b00000001110111001110001010111010;
   assign mem[245471:245440] = 32'b00000001100111011100010011010000;
   assign mem[245503:245472] = 32'b00000001111111010000011010010010;
   assign mem[245535:245504] = 32'b11111100110110100001011001101000;
   assign mem[245567:245536] = 32'b11110010010000000000111010100000;
   assign mem[245599:245568] = 32'b00000001011101000011010000011000;
   assign mem[245631:245600] = 32'b00000011100111010010101101011000;
   assign mem[245663:245632] = 32'b00000001100111011101100111100100;
   assign mem[245695:245664] = 32'b11111100010100010011011111000000;
   assign mem[245727:245696] = 32'b11111100001101101101010100111100;
   assign mem[245759:245728] = 32'b00000100100000001111111100100000;
   assign mem[245791:245760] = 32'b00001010001001000101010000000000;
   assign mem[245823:245792] = 32'b11110101100100011001010000010000;
   assign mem[245855:245824] = 32'b11111100001000101101000010011100;
   assign mem[245887:245856] = 32'b00000000010100111111010111100101;
   assign mem[245919:245888] = 32'b00000101010011010111001101000000;
   assign mem[245951:245920] = 32'b11111101101010110011100110000100;
   assign mem[245983:245952] = 32'b00000001010011011110101011111000;
   assign mem[246015:245984] = 32'b11111011011111110101011110111000;
   assign mem[246047:246016] = 32'b00000011101100010010000101001000;
   assign mem[246079:246048] = 32'b00000000000111100001011110111111;
   assign mem[246111:246080] = 32'b00001001000100101101011010110000;
   assign mem[246143:246112] = 32'b00000011101001111001100101010100;
   assign mem[246175:246144] = 32'b00000100110011001011001100101000;
   assign mem[246207:246176] = 32'b11110110000110000010010101000000;
   assign mem[246239:246208] = 32'b11111010001011010100100100101000;
   assign mem[246271:246240] = 32'b00000111000100010111100000010000;
   assign mem[246303:246272] = 32'b11111101011000101011111110000000;
   assign mem[246335:246304] = 32'b00001101000010011011111110010000;
   assign mem[246367:246336] = 32'b11111001110101111010100111001000;
   assign mem[246399:246368] = 32'b11101010110100011010111110100000;
   assign mem[246431:246400] = 32'b00000001101100111101110010111000;
   assign mem[246463:246432] = 32'b11111110101100100100110101101110;
   assign mem[246495:246464] = 32'b11111110100100100001110110000110;
   assign mem[246527:246496] = 32'b00000000010110010001010001100111;
   assign mem[246559:246528] = 32'b00001001111001100010001000010000;
   assign mem[246591:246560] = 32'b00000000010110010011011111101010;
   assign mem[246623:246592] = 32'b11111101001011101001001010001000;
   assign mem[246655:246624] = 32'b11110011110111110110101111100000;
   assign mem[246687:246656] = 32'b00000010111110001000111111111000;
   assign mem[246719:246688] = 32'b11111111000001111100110010100110;
   assign mem[246751:246720] = 32'b11110100010100001111000000010000;
   assign mem[246783:246752] = 32'b11110000000000110000101111100000;
   assign mem[246815:246784] = 32'b11111111101100101000010000110100;
   assign mem[246847:246816] = 32'b11111111111111000101001001001000;
   assign mem[246879:246848] = 32'b11111110010001101110011110010010;
   assign mem[246911:246880] = 32'b00000001111000100011100001110000;
   assign mem[246943:246912] = 32'b11110101011100001111110000110000;
   assign mem[246975:246944] = 32'b00000000000101110101001010000100;
   assign mem[247007:246976] = 32'b11111001111011011101101110101000;
   assign mem[247039:247008] = 32'b00000111011110001101111111001000;
   assign mem[247071:247040] = 32'b11111101011110011111100000101100;
   assign mem[247103:247072] = 32'b00000010000010100010100011001000;
   assign mem[247135:247104] = 32'b00000100000001001111011111011000;
   assign mem[247167:247136] = 32'b00000001101110101010001101110010;
   assign mem[247199:247168] = 32'b11111101100001110101110001010000;
   assign mem[247231:247200] = 32'b00000010010100010001101001001000;
   assign mem[247263:247232] = 32'b11111101000100001110100111110100;
   assign mem[247295:247264] = 32'b00000011001010001001011111011100;
   assign mem[247327:247296] = 32'b11110001011111001100001101110000;
   assign mem[247359:247328] = 32'b11111100100100110100010010010000;
   assign mem[247391:247360] = 32'b11111110111010011100011001101010;
   assign mem[247423:247392] = 32'b11111110100110101000000001010110;
   assign mem[247455:247424] = 32'b11111010011000111101101001111000;
   assign mem[247487:247456] = 32'b11111101011010111001110100011000;
   assign mem[247519:247488] = 32'b00000011011001000111100110110100;
   assign mem[247551:247520] = 32'b00000000010101000000111001010011;
   assign mem[247583:247552] = 32'b00000100011100100101101101100000;
   assign mem[247615:247584] = 32'b00000000101001010100110101011000;
   assign mem[247647:247616] = 32'b00000001010001010001000000111100;
   assign mem[247679:247648] = 32'b11111110010110101111000111010110;
   assign mem[247711:247680] = 32'b00000011110001011110111100101000;
   assign mem[247743:247712] = 32'b00000001011001110110110001001000;
   assign mem[247775:247744] = 32'b11111011111101111111000011100000;
   assign mem[247807:247776] = 32'b11110111010100110010110011010000;
   assign mem[247839:247808] = 32'b00000000001000001011010000000101;
   assign mem[247871:247840] = 32'b00000001101001000100110111000110;
   assign mem[247903:247872] = 32'b11111101111000011111010111011100;
   assign mem[247935:247904] = 32'b00001111000000000100111110000000;
   assign mem[247967:247936] = 32'b11110011010010110100110110100000;
   assign mem[247999:247968] = 32'b11111011110001110111001000101000;
   assign mem[248031:248000] = 32'b00000100001000101110101000110000;
   assign mem[248063:248032] = 32'b00000110100011100110001010000000;
   assign mem[248095:248064] = 32'b11111101001001100111010100000000;
   assign mem[248127:248096] = 32'b00000000110110010110010010010001;
   assign mem[248159:248128] = 32'b11111101110101010000000011110000;
   assign mem[248191:248160] = 32'b00000000100101111010000000001010;
   assign mem[248223:248192] = 32'b00000101101100010100110010100000;
   assign mem[248255:248224] = 32'b00000100110001010000101101001000;
   assign mem[248287:248256] = 32'b00000000011001111011100010001100;
   assign mem[248319:248288] = 32'b11111101100101111011100000100000;
   assign mem[248351:248320] = 32'b11111111110101111011101010111011;
   assign mem[248383:248352] = 32'b11110001010100110001111011100000;
   assign mem[248415:248384] = 32'b00000111011100001011000101101000;
   assign mem[248447:248416] = 32'b11111111110100010000100011010100;
   assign mem[248479:248448] = 32'b11111100011001001100101000110100;
   assign mem[248511:248480] = 32'b00000011110111100101001001100100;
   assign mem[248543:248512] = 32'b11111001110111000001010011100000;
   assign mem[248575:248544] = 32'b00001000010110010110101000110000;
   assign mem[248607:248576] = 32'b11110110010101110001110110000000;
   assign mem[248639:248608] = 32'b11110111101101111011011111100000;
   assign mem[248671:248640] = 32'b11110010000101111111100000010000;
   assign mem[248703:248672] = 32'b00000100111011100110001101010000;
   assign mem[248735:248704] = 32'b00000100010100111001101100010000;
   assign mem[248767:248736] = 32'b11111011011111010011011111000000;
   assign mem[248799:248768] = 32'b11110001110001111011111100010000;
   assign mem[248831:248800] = 32'b00000100100100101011110101000000;
   assign mem[248863:248832] = 32'b11111111000011100100000001101101;
   assign mem[248895:248864] = 32'b00001010000110110111001111100000;
   assign mem[248927:248896] = 32'b11111101000100001110001011001100;
   assign mem[248959:248928] = 32'b11111011101111110110100010101000;
   assign mem[248991:248960] = 32'b11110010000101101111010011100000;
   assign mem[249023:248992] = 32'b00000111010110010001001101101000;
   assign mem[249055:249024] = 32'b00000101101001101101000010100000;
   assign mem[249087:249056] = 32'b00000011001000010100111101110000;
   assign mem[249119:249088] = 32'b00000001110010000101010100100110;
   assign mem[249151:249120] = 32'b00000011111001111010100111000000;
   assign mem[249183:249152] = 32'b00000010010010011101001101011000;
   assign mem[249215:249184] = 32'b11111110001101011001111011111110;
   assign mem[249247:249216] = 32'b11111101001001010101010010110000;
   assign mem[249279:249248] = 32'b00000100010110000001100100010000;
   assign mem[249311:249280] = 32'b11111100001001101101110100111000;
   assign mem[249343:249312] = 32'b11111111100111111101100100001001;
   assign mem[249375:249344] = 32'b11110101111111001100010110010000;
   assign mem[249407:249376] = 32'b00000101000000000110101100111000;
   assign mem[249439:249408] = 32'b00000100010011101111110100001000;
   assign mem[249471:249440] = 32'b00000101000101001001100111000000;
   assign mem[249503:249472] = 32'b11110100010110010111110000110000;
   assign mem[249535:249504] = 32'b11111010011111110000110110101000;
   assign mem[249567:249536] = 32'b00000011010100111001000000111100;
   assign mem[249599:249568] = 32'b00000010011111001000101001111100;
   assign mem[249631:249600] = 32'b11111010000111010111110010101000;
   assign mem[249663:249632] = 32'b11100101001011011100100100100000;
   assign mem[249695:249664] = 32'b00000101101000101100010000110000;
   assign mem[249727:249696] = 32'b11111101001111000100100110001100;
   assign mem[249759:249728] = 32'b00001001100110110110010100010000;
   assign mem[249791:249760] = 32'b00000010010011001110110010111000;
   assign mem[249823:249792] = 32'b00001000000101011000001101100000;
   assign mem[249855:249824] = 32'b11101111110000100100110101000000;
   assign mem[249887:249856] = 32'b00000001001000000011100010010100;
   assign mem[249919:249888] = 32'b00000001010110011010010011111110;
   assign mem[249951:249920] = 32'b11111101010010111011100101010100;
   assign mem[249983:249952] = 32'b11110101100100101100111011100000;
   assign mem[250015:249984] = 32'b00001011110010101101111110110000;
   assign mem[250047:250016] = 32'b11111000010101110011110010001000;
   assign mem[250079:250048] = 32'b00001000111001011001001001110000;
   assign mem[250111:250080] = 32'b00001011010000001000110111010000;
   assign mem[250143:250112] = 32'b00001010111010111111000100110000;
   assign mem[250175:250144] = 32'b11110101101001110010010101000000;
   assign mem[250207:250176] = 32'b11111010001010111101000110111000;
   assign mem[250239:250208] = 32'b11110101101111000011001110010000;
   assign mem[250271:250240] = 32'b11111000001100001011111011101000;
   assign mem[250303:250272] = 32'b11110000001100001100111001000000;
   assign mem[250335:250304] = 32'b11111011101100110110001000010000;
   assign mem[250367:250336] = 32'b11111101010010011100000000110000;
   assign mem[250399:250368] = 32'b00000101110001011011111100011000;
   assign mem[250431:250400] = 32'b00000010010111000100101101101000;
   assign mem[250463:250432] = 32'b00000000101100001111110110110110;
   assign mem[250495:250464] = 32'b11101011000111110100101100000000;
   assign mem[250527:250496] = 32'b00000101011101111101000011100000;
   assign mem[250559:250528] = 32'b00000110110000111000011000111000;
   assign mem[250591:250560] = 32'b11110011001010110011100111100000;
   assign mem[250623:250592] = 32'b00000000100011000011010001100001;
   assign mem[250655:250624] = 32'b00000000000001010110111001010101;
   assign mem[250687:250656] = 32'b11111111110010011101111010010001;
   assign mem[250719:250688] = 32'b11110101110000011101100111000000;
   assign mem[250751:250720] = 32'b11111011001110000110111011010000;
   assign mem[250783:250752] = 32'b11111111001110100110100001111010;
   assign mem[250815:250784] = 32'b00000011001110101000100100000000;
   assign mem[250847:250816] = 32'b00000100101011100010000010100000;
   assign mem[250879:250848] = 32'b11111101100011010100110110100100;
   assign mem[250911:250880] = 32'b11110111011010000001111010110000;
   assign mem[250943:250912] = 32'b11101010100010111010000000100000;
   assign mem[250975:250944] = 32'b11110100110011111101111000000000;
   assign mem[251007:250976] = 32'b11111111011101111010110111100111;
   assign mem[251039:251008] = 32'b00000000101100010000001111110101;
   assign mem[251071:251040] = 32'b00000001100110111100101001111100;
   assign mem[251103:251072] = 32'b00000000111000000100011010110001;
   assign mem[251135:251104] = 32'b11111010111011011010111011001000;
   assign mem[251167:251136] = 32'b11111111110010100000100011010010;
   assign mem[251199:251168] = 32'b00001000001011010010001110010000;
   assign mem[251231:251200] = 32'b11110100101111111001010011000000;
   assign mem[251263:251232] = 32'b11111111011000011010100101111101;
   assign mem[251295:251264] = 32'b00000000010100101111100010000000;
   assign mem[251327:251296] = 32'b00000010110000011111111110011100;
   assign mem[251359:251328] = 32'b00000101101101001110111010011000;
   assign mem[251391:251360] = 32'b11111011100111100010011000001000;
   assign mem[251423:251392] = 32'b11110110001001011100000001010000;
   assign mem[251455:251424] = 32'b11111101000101101010011010111100;
   assign mem[251487:251456] = 32'b00000001110000111110000100100000;
   assign mem[251519:251488] = 32'b00000100011001110100111100111000;
   assign mem[251551:251520] = 32'b11111011110110101111011100100000;
   assign mem[251583:251552] = 32'b11111101011100101011101110000000;
   assign mem[251615:251584] = 32'b11111110001100100101101001000110;
   assign mem[251647:251616] = 32'b11111111011001110101101000100011;
   assign mem[251679:251648] = 32'b00001000101101011001100111010000;
   assign mem[251711:251680] = 32'b00001010011010111100000001100000;
   assign mem[251743:251712] = 32'b11111111100010001101111101101100;
   assign mem[251775:251744] = 32'b00000001111111000001101101111010;
   assign mem[251807:251776] = 32'b11111001010110000001000111011000;
   assign mem[251839:251808] = 32'b11111110001101100111111101111100;
   assign mem[251871:251840] = 32'b11101111010110111100101100100000;
   assign mem[251903:251872] = 32'b11101111101010111010111100000000;
   assign mem[251935:251904] = 32'b00000100011101000010101010000000;
   assign mem[251967:251936] = 32'b00001001110111011101000101110000;
   assign mem[251999:251968] = 32'b11111101010111001111111010001000;
   assign mem[252031:252000] = 32'b00000000001001000000101100100011;
   assign mem[252063:252032] = 32'b11111011010110000101111011001000;
   assign mem[252095:252064] = 32'b00000000101001000011011001110100;
   assign mem[252127:252096] = 32'b00000101101110110010010001100000;
   assign mem[252159:252128] = 32'b00000101010100111101100101000000;
   assign mem[252191:252160] = 32'b11111000010000010000011101101000;
   assign mem[252223:252192] = 32'b00000101101100011111101011100000;
   assign mem[252255:252224] = 32'b11111011101010110001011000010000;
   assign mem[252287:252256] = 32'b11111110001101110000111010110010;
   assign mem[252319:252288] = 32'b11111111000110100100011110001001;
   assign mem[252351:252320] = 32'b00000000000110000100011111000110;
   assign mem[252383:252352] = 32'b11111111110010110011000101111011;
   assign mem[252415:252384] = 32'b00001001000111110101101000000000;
   assign mem[252447:252416] = 32'b11111110100101011111110111100010;
   assign mem[252479:252448] = 32'b00000000100000010011001000101101;
   assign mem[252511:252480] = 32'b11110101101110101010010001000000;
   assign mem[252543:252512] = 32'b11111011100110110010111001000000;
   assign mem[252575:252544] = 32'b00000011110100011010010010111100;
   assign mem[252607:252576] = 32'b00000011001000111111101000100100;
   assign mem[252639:252608] = 32'b00000001010101110001101001001010;
   assign mem[252671:252640] = 32'b00000010010110100111000011010100;
   assign mem[252703:252672] = 32'b00000000111010101000000111101110;
   assign mem[252735:252704] = 32'b11110111000110101010110110100000;
   assign mem[252767:252736] = 32'b00000101001111100110010110101000;
   assign mem[252799:252768] = 32'b00000110111101110110101100110000;
   assign mem[252831:252800] = 32'b00000011011101101001001111110100;
   assign mem[252863:252832] = 32'b00000010110100011110110111100100;
   assign mem[252895:252864] = 32'b11111110100000010010101111000010;
   assign mem[252927:252896] = 32'b00000001100111000110111101010100;
   assign mem[252959:252928] = 32'b00000001100111010000110100011000;
   assign mem[252991:252960] = 32'b11111100101100100101011000000100;
   assign mem[253023:252992] = 32'b00000101010000111011110100101000;
   assign mem[253055:253024] = 32'b11111000001101110000010110001000;
   assign mem[253087:253056] = 32'b00000001011001100110000101101110;
   assign mem[253119:253088] = 32'b11111111101011011011111001000101;
   assign mem[253151:253120] = 32'b11111100011100111111000001011100;
   assign mem[253183:253152] = 32'b00000011101100111110000111011100;
   assign mem[253215:253184] = 32'b11110010111101011000001101010000;
   assign mem[253247:253216] = 32'b00000101000011110010101101011000;
   assign mem[253279:253248] = 32'b11111011001000101111111100111000;
   assign mem[253311:253280] = 32'b00000001110111110111101001110100;
   assign mem[253343:253312] = 32'b11111100101010111100111010001100;
   assign mem[253375:253344] = 32'b11111010000001011101110100111000;
   assign mem[253407:253376] = 32'b00001000100011100010110010110000;
   assign mem[253439:253408] = 32'b11111111011000100011010100110011;
   assign mem[253471:253440] = 32'b11111110000010000101100001011100;
   assign mem[253503:253472] = 32'b00000000001011110111100011111010;
   assign mem[253535:253504] = 32'b11110110010010100001000100110000;
   assign mem[253567:253536] = 32'b00000000000110011000011110001001;
   assign mem[253599:253568] = 32'b11111110101001011100100111000100;
   assign mem[253631:253600] = 32'b00000100011110011010110101111000;
   assign mem[253663:253632] = 32'b11110101110100000011001100000000;
   assign mem[253695:253664] = 32'b11111001100011110000010001010000;
   assign mem[253727:253696] = 32'b00001011011010010000011100010000;
   assign mem[253759:253728] = 32'b00000000101010111011000010111011;
   assign mem[253791:253760] = 32'b00000001000111001010010111010010;
   assign mem[253823:253792] = 32'b00000111100001100101000011111000;
   assign mem[253855:253824] = 32'b11111101101011000101011110000100;
   assign mem[253887:253856] = 32'b11110000100010110001100111100000;
   assign mem[253919:253888] = 32'b11111100100111011010110001000000;
   assign mem[253951:253920] = 32'b00000101010011100110011100100000;
   assign mem[253983:253952] = 32'b00000000100101000001001011011001;
   assign mem[254015:253984] = 32'b00001100011101010001101000110000;
   assign mem[254047:254016] = 32'b11110111100110011000100100010000;
   assign mem[254079:254048] = 32'b11111011111011100111000011101000;
   assign mem[254111:254080] = 32'b00001001010001101011000001110000;
   assign mem[254143:254112] = 32'b11111010000100101100101110010000;
   assign mem[254175:254144] = 32'b11110101100000000011011001010000;
   assign mem[254207:254176] = 32'b11101110011001110100101101100000;
   assign mem[254239:254208] = 32'b00000100111001100011111011011000;
   assign mem[254271:254240] = 32'b00000001011000100101001100101110;
   assign mem[254303:254272] = 32'b00000001011001000010100110101000;
   assign mem[254335:254304] = 32'b00000110011011110101100101001000;
   assign mem[254367:254336] = 32'b00000110110011100100100100110000;
   assign mem[254399:254368] = 32'b11111111011000110101101001110000;
   assign mem[254431:254400] = 32'b11110001011110111010100000110000;
   assign mem[254463:254432] = 32'b00001001111010111101000110100000;
   assign mem[254495:254464] = 32'b00000100000010101001100011010000;
   assign mem[254527:254496] = 32'b00000000000000100111110100111010;
   assign mem[254559:254528] = 32'b11111000000101111000101101000000;
   assign mem[254591:254560] = 32'b11111010001001100100000010110000;
   assign mem[254623:254592] = 32'b00001010001101110111001001100000;
   assign mem[254655:254624] = 32'b00000111000101000111010011011000;
   assign mem[254687:254656] = 32'b11111010100000100111001101011000;
   assign mem[254719:254688] = 32'b11111100010001110111000001110100;
   assign mem[254751:254720] = 32'b11110100001000100110001001100000;
   assign mem[254783:254752] = 32'b11101011100011110100010111000000;
   assign mem[254815:254784] = 32'b11111101111010010011111001000100;
   assign mem[254847:254816] = 32'b00000000000111111000101100001001;
   assign mem[254879:254848] = 32'b00001001110011100111011000110000;
   assign mem[254911:254880] = 32'b00000100000111101100100011101000;
   assign mem[254943:254912] = 32'b00000000101010101110010101010101;
   assign mem[254975:254944] = 32'b11110001111011111101101010110000;
   assign mem[255007:254976] = 32'b00000001101011111101111111011100;
   assign mem[255039:255008] = 32'b00000110001111100110000100001000;
   assign mem[255071:255040] = 32'b11101100110001101000001000000000;
   assign mem[255103:255072] = 32'b00000000100101100011010001010101;
   assign mem[255135:255104] = 32'b00000111111001000100010001111000;
   assign mem[255167:255136] = 32'b00000010101111000100111000101100;
   assign mem[255199:255168] = 32'b00000110001010111000011100101000;
   assign mem[255231:255200] = 32'b00000101110101110001100100111000;
   assign mem[255263:255232] = 32'b00000101010111101010010011100000;
   assign mem[255295:255264] = 32'b00001000100110001100110000010000;
   assign mem[255327:255296] = 32'b11111000111011110110100001000000;
   assign mem[255359:255328] = 32'b11110111111100100011000101110000;
   assign mem[255391:255360] = 32'b00000100100001111001111010110000;
   assign mem[255423:255392] = 32'b00001000001100111011001110010000;
   assign mem[255455:255424] = 32'b11111110101001101111111101001100;
   assign mem[255487:255456] = 32'b11111001011011110011101111000000;
   assign mem[255519:255488] = 32'b11111011000111010111001101111000;
   assign mem[255551:255520] = 32'b00000101110001011100000101100000;
   assign mem[255583:255552] = 32'b11111111111111111111010111011011;
   assign mem[255615:255584] = 32'b00000010000101100000011111101000;
   assign mem[255647:255616] = 32'b11111111110010111101100001010010;
   assign mem[255679:255648] = 32'b11110111010000110000000110000000;
   assign mem[255711:255680] = 32'b00000010001000001101111010011000;
   assign mem[255743:255712] = 32'b11101111001010100100011011000000;
   assign mem[255775:255744] = 32'b11110110101010010110000111110000;
   assign mem[255807:255776] = 32'b11111110010111000100010000110100;
   assign mem[255839:255808] = 32'b00000010000100001011001110001000;
   assign mem[255871:255840] = 32'b00000011100101001010110101011000;
   assign mem[255903:255872] = 32'b11111111011001010001110000001110;
   assign mem[255935:255904] = 32'b00000010011001010000011101100000;
   assign mem[255967:255936] = 32'b11111010111101000011011001011000;
   assign mem[255999:255968] = 32'b00000111010001110000001100011000;
   assign mem[256031:256000] = 32'b00000000010100101001100100100111;
   assign mem[256063:256032] = 32'b11111110110011011000100101100110;
   assign mem[256095:256064] = 32'b00000000110100100010011011110001;
   assign mem[256127:256096] = 32'b00000010010000100010011100110000;
   assign mem[256159:256128] = 32'b11111100001001001101100101100000;
   assign mem[256191:256160] = 32'b11111101111001111001010001001000;
   assign mem[256223:256192] = 32'b00000000101000111100010010101010;
   assign mem[256255:256224] = 32'b11111111010001000110001001010110;
   assign mem[256287:256256] = 32'b00000000100101011110111111111100;
   assign mem[256319:256288] = 32'b11111100101100110010010001010100;
   assign mem[256351:256320] = 32'b00000101001111001101100010100000;
   assign mem[256383:256352] = 32'b00000011110001010001000011111000;
   assign mem[256415:256384] = 32'b00000000011101110100100001110100;
   assign mem[256447:256416] = 32'b00000010100111000110100111011100;
   assign mem[256479:256448] = 32'b11111100111110111000101110001000;
   assign mem[256511:256480] = 32'b00000000100100011001100011100000;
   assign mem[256543:256512] = 32'b00000110011110101011001001001000;
   assign mem[256575:256544] = 32'b00000011000101100011001000111100;
   assign mem[256607:256576] = 32'b11111010100110000011100010110000;
   assign mem[256639:256608] = 32'b11111000001101010011111000100000;
   assign mem[256671:256640] = 32'b11111110100100110111010001010100;
   assign mem[256703:256672] = 32'b11111011001000110110011101110000;
   assign mem[256735:256704] = 32'b11111101010001101110101011101100;
   assign mem[256767:256736] = 32'b11111100110011111010001010001000;
   assign mem[256799:256768] = 32'b00000111001011110100001110110000;
   assign mem[256831:256800] = 32'b00000010111101011000000011000100;
   assign mem[256863:256832] = 32'b00000010100011100010110111011100;
   assign mem[256895:256864] = 32'b11111011011110011101100110000000;
   assign mem[256927:256896] = 32'b11111100001000010000000011010100;
   assign mem[256959:256928] = 32'b00000010100100100000101110101100;
   assign mem[256991:256960] = 32'b00000100011111101001110100111000;
   assign mem[257023:256992] = 32'b00000010100100011000111110110000;
   assign mem[257055:257024] = 32'b11111011100011100000101010001000;
   assign mem[257087:257056] = 32'b00001010101010101000001111100000;
   assign mem[257119:257088] = 32'b11111111101111111001100001111010;
   assign mem[257151:257120] = 32'b11111110101011010010010000001010;
   assign mem[257183:257152] = 32'b11111111010001000011010010100101;
   assign mem[257215:257184] = 32'b00010010010011110110110101100000;
   assign mem[257247:257216] = 32'b11100110000111100001000000000000;
   assign mem[257279:257248] = 32'b11111011000010010000000010110000;
   assign mem[257311:257280] = 32'b11111010100101000011100100111000;
   assign mem[257343:257312] = 32'b11100100000011111100011110100000;
   assign mem[257375:257344] = 32'b00000110111101111110001011111000;
   assign mem[257407:257376] = 32'b11111101011011000101110101101100;
   assign mem[257439:257408] = 32'b00000101001000111011000000111000;
   assign mem[257471:257440] = 32'b00000100001010111000110011100000;
   assign mem[257503:257472] = 32'b11111110011111101110110100010000;
   assign mem[257535:257504] = 32'b11111100011100111110101000100000;
   assign mem[257567:257536] = 32'b00000000001101111110111101101010;
   assign mem[257599:257568] = 32'b11111011011001001011110111111000;
   assign mem[257631:257600] = 32'b11110110011110101100000001110000;
   assign mem[257663:257632] = 32'b00000011001110000011000101001000;
   assign mem[257695:257664] = 32'b00000100011000000100010110001000;
   assign mem[257727:257696] = 32'b11111100011110111111001101011000;
   assign mem[257759:257728] = 32'b00000011101100110100111000001100;
   assign mem[257791:257760] = 32'b00000100110000011010110001101000;
   assign mem[257823:257792] = 32'b00000001100011101100011011111110;
   assign mem[257855:257824] = 32'b11110101000111010011010000010000;
   assign mem[257887:257856] = 32'b00000001110100011001111011000000;
   assign mem[257919:257888] = 32'b11111110000100010000111101100000;
   assign mem[257951:257920] = 32'b11111100111011111100110011110000;
   assign mem[257983:257952] = 32'b11110110111001110010101101100000;
   assign mem[258015:257984] = 32'b11110011101111011000101101000000;
   assign mem[258047:258016] = 32'b11111101110100100000011000100000;
   assign mem[258079:258048] = 32'b00000110100011001011001010011000;
   assign mem[258111:258080] = 32'b00000011110101011100001000000100;
   assign mem[258143:258112] = 32'b00000001011110000110110100011110;
   assign mem[258175:258144] = 32'b11110000010100011010100000100000;
   assign mem[258207:258176] = 32'b00000101000000000001001011011000;
   assign mem[258239:258208] = 32'b00000110011010000101011110010000;
   assign mem[258271:258240] = 32'b11111010101000000001100100000000;
   assign mem[258303:258272] = 32'b00000000010000101110110010001101;
   assign mem[258335:258304] = 32'b00000101110100101000111000100000;
   assign mem[258367:258336] = 32'b00000111110011000100110110100000;
   assign mem[258399:258368] = 32'b11110011011011110100101001100000;
   assign mem[258431:258400] = 32'b11110111111001000101110100000000;
   assign mem[258463:258432] = 32'b11111000010111011101011111001000;
   assign mem[258495:258464] = 32'b00000110011000101000010001001000;
   assign mem[258527:258496] = 32'b11101111110000111111111111100000;
   assign mem[258559:258528] = 32'b00000000110001110001110001000011;
   assign mem[258591:258560] = 32'b00001001001001100100011101000000;
   assign mem[258623:258592] = 32'b00000101010110010000101101011000;
   assign mem[258655:258624] = 32'b11111001001001000000000000111000;
   assign mem[258687:258656] = 32'b11111001001001011101010110111000;
   assign mem[258719:258688] = 32'b00000100101000010110000111000000;
   assign mem[258751:258720] = 32'b11111011110011011111000010100000;
   assign mem[258783:258752] = 32'b11110111010010100010010000100000;
   assign mem[258815:258784] = 32'b11111110010000000101111101110100;
   assign mem[258847:258816] = 32'b00000101010110000000101100010000;
   assign mem[258879:258848] = 32'b11111110110111100111011000000010;
   assign mem[258911:258880] = 32'b11111111110100001011111101111000;
   assign mem[258943:258912] = 32'b11110110111101001101000101000000;
   assign mem[258975:258944] = 32'b00000010100100111011101100101000;
   assign mem[259007:258976] = 32'b00000100111010101001101111010000;
   assign mem[259039:259008] = 32'b11111101111110011110101001110000;
   assign mem[259071:259040] = 32'b00000001100100101001100000001010;
   assign mem[259103:259072] = 32'b00000001000101010010011100111100;
   assign mem[259135:259104] = 32'b00000010100011011011111110101100;
   assign mem[259167:259136] = 32'b11111001101110100010110001111000;
   assign mem[259199:259168] = 32'b11111101101000110001010101110000;
   assign mem[259231:259200] = 32'b00000001110100101100101011011110;
   assign mem[259263:259232] = 32'b11110101111111011001001100010000;
   assign mem[259295:259264] = 32'b00001000000011110010100110010000;
   assign mem[259327:259296] = 32'b00001000000110110110110110010000;
   assign mem[259359:259328] = 32'b11111100100100001011111100100100;
   assign mem[259391:259360] = 32'b00000100010101111100101011110000;
   assign mem[259423:259392] = 32'b11101011100000001001010010100000;
   assign mem[259455:259424] = 32'b11111101100010101011111101000000;
   assign mem[259487:259456] = 32'b11101011000100001101001101100000;
   assign mem[259519:259488] = 32'b00000110100001001111111101111000;
   assign mem[259551:259520] = 32'b00001011011001111010011000010000;
   assign mem[259583:259552] = 32'b00000100110111100011110110000000;
   assign mem[259615:259584] = 32'b11111101101010000101110100111000;
   assign mem[259647:259616] = 32'b11101111001001001010000101000000;
   assign mem[259679:259648] = 32'b00000000100000111111001101011101;
   assign mem[259711:259680] = 32'b00001000001101111111011100110000;
   assign mem[259743:259712] = 32'b11111110010011010110010101110100;
   assign mem[259775:259744] = 32'b11111011110000011110000000110000;
   assign mem[259807:259776] = 32'b00000001010100111100111110110000;
   assign mem[259839:259808] = 32'b11110100000011001101101001010000;
   assign mem[259871:259840] = 32'b11111110100110111000001101101110;
   assign mem[259903:259872] = 32'b11111010110000110100011001110000;
   assign mem[259935:259904] = 32'b11111001101010111101111101111000;
   assign mem[259967:259936] = 32'b00000001000100110011011111010000;
   assign mem[259999:259968] = 32'b00000100011010001100111101011000;
   assign mem[260031:260000] = 32'b00000010101101011100011000110100;
   assign mem[260063:260032] = 32'b00000010101100100000110010011100;
   assign mem[260095:260064] = 32'b11101101111100111011110101000000;
   assign mem[260127:260096] = 32'b00000001100011110111101010110010;
   assign mem[260159:260128] = 32'b00001000011111110001001001000000;
   assign mem[260191:260160] = 32'b11101101101000010000101011100000;
   assign mem[260223:260192] = 32'b00001001011010111011100100110000;
   assign mem[260255:260224] = 32'b00000101101110001101101010011000;
   assign mem[260287:260256] = 32'b11110011011101010111111100000000;
   assign mem[260319:260288] = 32'b11111100010000100110101110011000;
   assign mem[260351:260320] = 32'b00000011010010011100011000000100;
   assign mem[260383:260352] = 32'b11110111000011000101011110100000;
   assign mem[260415:260384] = 32'b11111000101111100101111111000000;
   assign mem[260447:260416] = 32'b00001101000010010101110000000000;
   assign mem[260479:260448] = 32'b11111100111100100111010111100000;
   assign mem[260511:260480] = 32'b11111101110000100001100111001100;
   assign mem[260543:260512] = 32'b00000010011000100110011010101000;
   assign mem[260575:260544] = 32'b11111101110111000001111011000100;
   assign mem[260607:260576] = 32'b11111011100101110101001000110000;
   assign mem[260639:260608] = 32'b00000011000011001101010000011000;
   assign mem[260671:260640] = 32'b00000000100111000001111101111010;
   assign mem[260703:260672] = 32'b11110111100110111111001101110000;
   assign mem[260735:260704] = 32'b11111111101000000011000011011011;
   assign mem[260767:260736] = 32'b11111101111101110101110011010100;
   assign mem[260799:260768] = 32'b00000100001011110010101001101000;
   assign mem[260831:260800] = 32'b00000011010011101111111111110000;
   assign mem[260863:260832] = 32'b11111111011110101001001010101111;
   assign mem[260895:260864] = 32'b00000011000111100011110101111100;
   assign mem[260927:260896] = 32'b00000000001010111110001011011000;
   assign mem[260959:260928] = 32'b00000010111010000111000110111100;
   assign mem[260991:260960] = 32'b11111111010010001001101101001110;
   assign mem[261023:260992] = 32'b00000011000101110000111111111100;
   assign mem[261055:261024] = 32'b11111110110000000001011100111000;
   assign mem[261087:261056] = 32'b11111011110001100101000111010000;
   assign mem[261119:261088] = 32'b11111101010110001100110011001100;
   assign mem[261151:261120] = 32'b00000010101000010010001011000100;
   assign mem[261183:261152] = 32'b00000001001110011110001111011100;
   assign mem[261215:261184] = 32'b11111000100011001111110000010000;
   assign mem[261247:261216] = 32'b11111101101011110001110011100000;
   assign mem[261279:261248] = 32'b00000000111111111110000100000010;
   assign mem[261311:261280] = 32'b00000011111111110100101000101100;
   assign mem[261343:261312] = 32'b00000001110111100100110011101100;
   assign mem[261375:261344] = 32'b00000010100111100101101111110000;
   assign mem[261407:261376] = 32'b00000010100000101011110110001100;
   assign mem[261439:261408] = 32'b11111100001111111110000101010000;
   assign mem[261471:261440] = 32'b11111001000001111100010010110000;
   assign mem[261503:261472] = 32'b00000101010010001111000110000000;
   assign mem[261535:261504] = 32'b00000000011000101110100110000011;
   assign mem[261567:261536] = 32'b00000111000000110000110000101000;
   assign mem[261599:261568] = 32'b11110011100010110001111000000000;
   assign mem[261631:261600] = 32'b00000010110010101110110010010100;
   assign mem[261663:261632] = 32'b00000101101101100100011111010000;
   assign mem[261695:261664] = 32'b00000110001000110000001110011000;
   assign mem[261727:261696] = 32'b11111011011000010110010000011000;
   assign mem[261759:261728] = 32'b11111010001111111000001110000000;
   assign mem[261791:261760] = 32'b11111100011010010111000100011000;
   assign mem[261823:261792] = 32'b11111010111010101000010011011000;
   assign mem[261855:261824] = 32'b00000000111001000111110100011001;
   assign mem[261887:261856] = 32'b11111101010111111010000111000100;
   assign mem[261919:261888] = 32'b11111011101110111110100110101000;
   assign mem[261951:261920] = 32'b11111011001010000010011110000000;
   assign mem[261983:261952] = 32'b00000010011001111000010011110100;
   assign mem[262015:261984] = 32'b11111101001000111000001101101000;
   assign mem[262047:262016] = 32'b00000101011111011111001000110000;
   assign mem[262079:262048] = 32'b00000111011011000011010101100000;
   assign mem[262111:262080] = 32'b11111011011001111001111110101000;
   assign mem[262143:262112] = 32'b00000100100001010101101110000000;
   assign mem[262175:262144] = 32'b00000000111110010001011100100100;
   assign mem[262207:262176] = 32'b00000000110011110100111100111001;
   assign mem[262239:262208] = 32'b11111000101000111001111111000000;
   assign mem[262271:262240] = 32'b11111111001110100111001101100111;
   assign mem[262303:262272] = 32'b11111010101111100110100100100000;
   assign mem[262335:262304] = 32'b00000110101111001010110111100000;
   assign mem[262367:262336] = 32'b11111101101111001000001111110000;
   assign mem[262399:262368] = 32'b11111000100111101110001010111000;
   assign mem[262431:262400] = 32'b11111001001000100010010010100000;
   assign mem[262463:262432] = 32'b11110100011011101110110111100000;
   assign mem[262495:262464] = 32'b11110111101111011010010000010000;
   assign mem[262527:262496] = 32'b00000011011110111000000001111000;
   assign mem[262559:262528] = 32'b00001000101010100010010010000000;
   assign mem[262591:262560] = 32'b11111110011010111011111011100110;
   assign mem[262623:262592] = 32'b11111100011010001001001000000000;
   assign mem[262655:262624] = 32'b00000000010100101010000000111110;
   assign mem[262687:262656] = 32'b11111110000010111100110010100000;
   assign mem[262719:262688] = 32'b00000111111010110100010111101000;
   assign mem[262751:262720] = 32'b11110100001100000001000001110000;
   assign mem[262783:262752] = 32'b11101111100111010110001101100000;
   assign mem[262815:262784] = 32'b00000000101101011101001010110011;
   assign mem[262847:262816] = 32'b00000011001110010011110001001100;
   assign mem[262879:262848] = 32'b00000111010010001010011111010000;
   assign mem[262911:262880] = 32'b00000010111111010101101010111000;
   assign mem[262943:262912] = 32'b00000100010011111001101000011000;
   assign mem[262975:262944] = 32'b11110101000110101101000011000000;
   assign mem[263007:262976] = 32'b11111111101111011101111111000001;
   assign mem[263039:263008] = 32'b00000001010000111110010011101100;
   assign mem[263071:263040] = 32'b11111101100110100110001101010000;
   assign mem[263103:263072] = 32'b00000001101110111001010000010110;
   assign mem[263135:263104] = 32'b11111010000101000100010100101000;
   assign mem[263167:263136] = 32'b00000110010101100010101011101000;
   assign mem[263199:263168] = 32'b11111110111111111110101000100000;
   assign mem[263231:263200] = 32'b00000011001100000001000001100100;
   assign mem[263263:263232] = 32'b11111110100000101010110000010010;
   assign mem[263295:263264] = 32'b00000010011001110100010111010100;
   assign mem[263327:263296] = 32'b11111100010001111010100110001000;
   assign mem[263359:263328] = 32'b11111110001000100111100010100010;
   assign mem[263391:263360] = 32'b00000100000111001100110111000000;
   assign mem[263423:263392] = 32'b00000001101000000010110000001010;
   assign mem[263455:263424] = 32'b11110101110111010011011111000000;
   assign mem[263487:263456] = 32'b11111001101000010001011010110000;
   assign mem[263519:263488] = 32'b00000011010010100100101011000000;
   assign mem[263551:263520] = 32'b11111110111000111001001000100000;
   assign mem[263583:263552] = 32'b00000000111000010011101110001111;
   assign mem[263615:263584] = 32'b00000101100111001111110101011000;
   assign mem[263647:263616] = 32'b11110011111101100110010000100000;
   assign mem[263679:263648] = 32'b00000100001110010101001011110000;
   assign mem[263711:263680] = 32'b00000110111001101000110101111000;
   assign mem[263743:263712] = 32'b00001010010110011010011111100000;
   assign mem[263775:263744] = 32'b11111011101100100000010100110000;
   assign mem[263807:263776] = 32'b00000100001000000010011111011000;
   assign mem[263839:263808] = 32'b11111010110111010100100010111000;
   assign mem[263871:263840] = 32'b11111110010100111110101111100000;
   assign mem[263903:263872] = 32'b11111001101101000101111100011000;
   assign mem[263935:263904] = 32'b11111001101010110101100001101000;
   assign mem[263967:263936] = 32'b11111011010011001100101010111000;
   assign mem[263999:263968] = 32'b00000000010010010001110101111100;
   assign mem[264031:264000] = 32'b11111101101101100010101000100100;
   assign mem[264063:264032] = 32'b11111010010000010100000110101000;
   assign mem[264095:264064] = 32'b11111100011000101001101000011100;
   assign mem[264127:264096] = 32'b11111100101010100111000010110000;
   assign mem[264159:264128] = 32'b00000010100100111011110011000100;
   assign mem[264191:264160] = 32'b00000000011001011111110111001001;
   assign mem[264223:264192] = 32'b11110001101010001001000110110000;
   assign mem[264255:264224] = 32'b11111100111101100110000001000100;
   assign mem[264287:264256] = 32'b00000111100010010111011100100000;
   assign mem[264319:264288] = 32'b00000100100110001101101010110000;
   assign mem[264351:264320] = 32'b11111010011001110100100001110000;
   assign mem[264383:264352] = 32'b11111000010001010010001010110000;
   assign mem[264415:264384] = 32'b00001100111010011001000010010000;
   assign mem[264447:264416] = 32'b11111010010111011110011000111000;
   assign mem[264479:264448] = 32'b11111011001111011110010001101000;
   assign mem[264511:264480] = 32'b00001000010111010101011011000000;
   assign mem[264543:264512] = 32'b00001001000110110101101011010000;
   assign mem[264575:264544] = 32'b00000011011101110010001100110100;
   assign mem[264607:264576] = 32'b11111001101110001111000110011000;
   assign mem[264639:264608] = 32'b11110110111000110111011011000000;
   assign mem[264671:264640] = 32'b11111011010100000101001000110000;
   assign mem[264703:264672] = 32'b00000010100010011101100111111000;
   assign mem[264735:264704] = 32'b00000100010100100110001001101000;
   assign mem[264767:264736] = 32'b11110110011110111010101010000000;
   assign mem[264799:264768] = 32'b11111100011100011100010111101100;
   assign mem[264831:264800] = 32'b00000001000011011100011101011100;
   assign mem[264863:264832] = 32'b00000001010111110000111111010000;
   assign mem[264895:264864] = 32'b11111010110101100001001011011000;
   assign mem[264927:264896] = 32'b00001101000000100010001101010000;
   assign mem[264959:264928] = 32'b11111010010010110011100000101000;
   assign mem[264991:264960] = 32'b11110100011001001010101100010000;
   assign mem[265023:264992] = 32'b00000000101001100011110101100000;
   assign mem[265055:265024] = 32'b00001000011011100011110010000000;
   assign mem[265087:265056] = 32'b00001000010000101110000000000000;
   assign mem[265119:265088] = 32'b11110111100010110000101011010000;
   assign mem[265151:265120] = 32'b11111110010110010001100011010000;
   assign mem[265183:265152] = 32'b00001010110000111010110011010000;
   assign mem[265215:265184] = 32'b00000011011110010011000000001000;
   assign mem[265247:265216] = 32'b11110110001100100010100101000000;
   assign mem[265279:265248] = 32'b11111110010100101111001100001100;
   assign mem[265311:265280] = 32'b00000001100100001001101110110100;
   assign mem[265343:265312] = 32'b00000100111001000010111100111000;
   assign mem[265375:265344] = 32'b00000000111110111011101100010010;
   assign mem[265407:265376] = 32'b00000011110010101010000110101100;
   assign mem[265439:265408] = 32'b11110110111100011110011000010000;
   assign mem[265471:265440] = 32'b00000001010010100011110111101010;
   assign mem[265503:265472] = 32'b00001000011000100110001010000000;
   assign mem[265535:265504] = 32'b00000000111101000111011001000010;
   assign mem[265567:265536] = 32'b11110110101100000111010111010000;
   assign mem[265599:265568] = 32'b11110111010011000100000110000000;
   assign mem[265631:265600] = 32'b11101010011111111100011100000000;
   assign mem[265663:265632] = 32'b00000110110010100100011011110000;
   assign mem[265695:265664] = 32'b11111000100110101001010011111000;
   assign mem[265727:265696] = 32'b00000010001111011101011111010100;
   assign mem[265759:265728] = 32'b11110101101000111100001001110000;
   assign mem[265791:265760] = 32'b00000110111110010010100010000000;
   assign mem[265823:265792] = 32'b00000000011010000010010001011110;
   assign mem[265855:265824] = 32'b00000110111110101010111000001000;
   assign mem[265887:265856] = 32'b11111111111110110101000100111110;
   assign mem[265919:265888] = 32'b11110111000110111011010010000000;
   assign mem[265951:265920] = 32'b11101110111001111010000110000000;
   assign mem[265983:265952] = 32'b00000011011110010001000000011100;
   assign mem[266015:265984] = 32'b00000000010100011001010111111010;
   assign mem[266047:266016] = 32'b11111000101010100011011111010000;
   assign mem[266079:266048] = 32'b11110001111100001001000111010000;
   assign mem[266111:266080] = 32'b00000001110001000100010111101100;
   assign mem[266143:266112] = 32'b11111111100100001010101001011001;
   assign mem[266175:266144] = 32'b00001000111010010111010110100000;
   assign mem[266207:266176] = 32'b00000010110101001011110001111100;
   assign mem[266239:266208] = 32'b11111001101001111111011011011000;
   assign mem[266271:266240] = 32'b00000000011001010110111001110101;
   assign mem[266303:266272] = 32'b11110110011011111011010111110000;
   assign mem[266335:266304] = 32'b11111111111100100100101101010111;
   assign mem[266367:266336] = 32'b00001011111111000000111000000000;
   assign mem[266399:266368] = 32'b11111101110001011001101001110100;
   assign mem[266431:266400] = 32'b11111010111100010001111001001000;
   assign mem[266463:266432] = 32'b00000111000010011101011100010000;
   assign mem[266495:266464] = 32'b00000100101111110110011010100000;
   assign mem[266527:266496] = 32'b00001000000101101111010100010000;
   assign mem[266559:266528] = 32'b11110101101001010011100101010000;
   assign mem[266591:266560] = 32'b00000011000010011111000010011000;
   assign mem[266623:266592] = 32'b00000100010011111110110001001000;
   assign mem[266655:266624] = 32'b00000010010111000010110100010000;
   assign mem[266687:266656] = 32'b00000010000010111000011001110000;
   assign mem[266719:266688] = 32'b11110100110110100111001101110000;
   assign mem[266751:266720] = 32'b00001000001101110111101100100000;
   assign mem[266783:266752] = 32'b00000111100101001111101001010000;
   assign mem[266815:266784] = 32'b11110110100110001000011010000000;
   assign mem[266847:266816] = 32'b11101100100101011110011110000000;
   assign mem[266879:266848] = 32'b00000101101011001000101100100000;
   assign mem[266911:266880] = 32'b11111110001101111101101110001110;
   assign mem[266943:266912] = 32'b11111111000010011111011011011011;
   assign mem[266975:266944] = 32'b11110111101001000011110011010000;
   assign mem[267007:266976] = 32'b00000100100101110100001110011000;
   assign mem[267039:267008] = 32'b11110110100010101101111001000000;
   assign mem[267071:267040] = 32'b00000101010000101000000010110000;
   assign mem[267103:267072] = 32'b00000101101100011111011100101000;
   assign mem[267135:267104] = 32'b11111110110101011011111010101110;
   assign mem[267167:267136] = 32'b00000000101010011011101011100111;
   assign mem[267199:267168] = 32'b11111110011110101111001101010100;
   assign mem[267231:267200] = 32'b00000010010011111001100101110100;
   assign mem[267263:267232] = 32'b11110111111000001000101000110000;
   assign mem[267295:267264] = 32'b11110101110111010111010111010000;
   assign mem[267327:267296] = 32'b00000111000101111101110100111000;
   assign mem[267359:267328] = 32'b11110000101111001110100010100000;
   assign mem[267391:267360] = 32'b00000110100111110111110110100000;
   assign mem[267423:267392] = 32'b11111010011111110101100000101000;
   assign mem[267455:267424] = 32'b00000010011111010001000101001100;
   assign mem[267487:267456] = 32'b00000000000010110100111011000011;
   assign mem[267519:267488] = 32'b00000010001101000111110101001100;
   assign mem[267551:267520] = 32'b11111110111010111000000100101010;
   assign mem[267583:267552] = 32'b11110011100010011000100101000000;
   assign mem[267615:267584] = 32'b11111110011101101111101001000010;
   assign mem[267647:267616] = 32'b11111010011011011111000110101000;
   assign mem[267679:267648] = 32'b11110010101010110000011110100000;
   assign mem[267711:267680] = 32'b00000100111001100011111100001000;
   assign mem[267743:267712] = 32'b11111001001001100100110100111000;
   assign mem[267775:267744] = 32'b00000001100001010011010001000100;
   assign mem[267807:267776] = 32'b11111100111011001001100011110000;
   assign mem[267839:267808] = 32'b00000101010000111000110101000000;
   assign mem[267871:267840] = 32'b11111100000111110101001110001100;
   assign mem[267903:267872] = 32'b00000100000001100011011011001000;
   assign mem[267935:267904] = 32'b00000110010110000110000110010000;
   assign mem[267967:267936] = 32'b00000001001101100100101000110010;
   assign mem[267999:267968] = 32'b11111111010111001100010001110100;
   assign mem[268031:268000] = 32'b11100111110100100011010010100000;
   assign mem[268063:268032] = 32'b11111010001010010000011000011000;
   assign mem[268095:268064] = 32'b00000100000011111000001110001000;
   assign mem[268127:268096] = 32'b00000010110111011100010000000100;
   assign mem[268159:268128] = 32'b11111001101011111010111000100000;
   assign mem[268191:268160] = 32'b00000001010001000010000001100100;
   assign mem[268223:268192] = 32'b00000000001101110000101100101011;
   assign mem[268255:268224] = 32'b11111111000111111011111000110011;
   assign mem[268287:268256] = 32'b11110110110001000010110110000000;
   assign mem[268319:268288] = 32'b11111001101001101111001000011000;
   assign mem[268351:268320] = 32'b00000100110100001100100010001000;
   assign mem[268383:268352] = 32'b11111110100011001000110110010110;
   assign mem[268415:268384] = 32'b00000011100001001011000111000100;
   assign mem[268447:268416] = 32'b11111110011010111110111000001010;
   assign mem[268479:268448] = 32'b00000111101111111010000000001000;
   assign mem[268511:268480] = 32'b11110101000001001110100110100000;
   assign mem[268543:268512] = 32'b11111111101100011100110101101001;
   assign mem[268575:268544] = 32'b00000101010100010111010101101000;
   assign mem[268607:268576] = 32'b00000110101010111110011001110000;
   assign mem[268639:268608] = 32'b11111110010111010001100101000010;
   assign mem[268671:268640] = 32'b11101101000010001110100000100000;
   assign mem[268703:268672] = 32'b11111010110100010011111011100000;
   assign mem[268735:268704] = 32'b00000100101111111000000010010000;
   assign mem[268767:268736] = 32'b00000001011000010011010000100000;
   assign mem[268799:268768] = 32'b11111111000110000011001011010101;
   assign mem[268831:268800] = 32'b11110011101101000011101111100000;
   assign mem[268863:268832] = 32'b11111110001010011101011111011100;
   assign mem[268895:268864] = 32'b00000101100001000101101011000000;
   assign mem[268927:268896] = 32'b11110111011111100001010011110000;
   assign mem[268959:268928] = 32'b11110101111100110010100111000000;
   assign mem[268991:268960] = 32'b00001000000000001000101001100000;
   assign mem[269023:268992] = 32'b00000111111101111100101000110000;
   assign mem[269055:269024] = 32'b11110001101110011001110111010000;
   assign mem[269087:269056] = 32'b11110011001011100011000101110000;
   assign mem[269119:269088] = 32'b00000100101001011010100001111000;
   assign mem[269151:269120] = 32'b00000010011111110001001101101100;
   assign mem[269183:269152] = 32'b11111011100101001000000010000000;
   assign mem[269215:269184] = 32'b00001000000001111001100110010000;
   assign mem[269247:269216] = 32'b11101010101000010000101110000000;
   assign mem[269279:269248] = 32'b00000010111100110011010100010100;
   assign mem[269311:269280] = 32'b00000111101111000111000111001000;
   assign mem[269343:269312] = 32'b11110101011101100110111110110000;
   assign mem[269375:269344] = 32'b00001001111000011000000101000000;
   assign mem[269407:269376] = 32'b11110001110110101001000111100000;
   assign mem[269439:269408] = 32'b11111010100010011111000111100000;
   assign mem[269471:269440] = 32'b11101011101111111101111011000000;
   assign mem[269503:269472] = 32'b11111010001000111111100000110000;
   assign mem[269535:269504] = 32'b11111001101011001101111001010000;
   assign mem[269567:269536] = 32'b00000010000101001001011000111100;
   assign mem[269599:269568] = 32'b00000011011010100111101110010100;
   assign mem[269631:269600] = 32'b00000001011110001100000000101010;
   assign mem[269663:269632] = 32'b00000101110110101010100110001000;
   assign mem[269695:269664] = 32'b00000110011110111011011000110000;
   assign mem[269727:269696] = 32'b00000101110110100001001010111000;
   assign mem[269759:269728] = 32'b00000010101001100100110101011000;
   assign mem[269791:269760] = 32'b00000101110000011001001110101000;
   assign mem[269823:269792] = 32'b11111111110111010000100000001101;
   assign mem[269855:269824] = 32'b11111100000100100010010100111000;
   assign mem[269887:269856] = 32'b00000000010001111011001011110011;
   assign mem[269919:269888] = 32'b11111011001111011100011111001000;
   assign mem[269951:269920] = 32'b11111110010111101111001011001000;
   assign mem[269983:269952] = 32'b00000000110001001000001110100000;
   assign mem[270015:269984] = 32'b00000100001001101101101011011000;
   assign mem[270047:270016] = 32'b00000000000110100010111010110100;
   assign mem[270079:270048] = 32'b00000000000110110011101110110000;
   assign mem[270111:270080] = 32'b11110100111111110001001111110000;
   assign mem[270143:270112] = 32'b11110011011101111011111101110000;
   assign mem[270175:270144] = 32'b00000101100011011100001110111000;
   assign mem[270207:270176] = 32'b00000011010110100000110000001100;
   assign mem[270239:270208] = 32'b00000110001100100011010101101000;
   assign mem[270271:270240] = 32'b00000001001100101010101110010010;
   assign mem[270303:270272] = 32'b00000100010010000111011110101000;
   assign mem[270335:270304] = 32'b00001011001110011111110100010000;
   assign mem[270367:270336] = 32'b00000010000101100001011010100000;
   assign mem[270399:270368] = 32'b11110000010000000100111111100000;
   assign mem[270431:270400] = 32'b11110000100111101000111100100000;
   assign mem[270463:270432] = 32'b11110111001001000010100000000000;
   assign mem[270495:270464] = 32'b11111101111010110100100011011100;
   assign mem[270527:270496] = 32'b00000011101010011100111100001000;
   assign mem[270559:270528] = 32'b11111000001010110010100101110000;
   assign mem[270591:270560] = 32'b00000100001101000011111101000000;
   assign mem[270623:270592] = 32'b00001000010010001101101010100000;
   assign mem[270655:270624] = 32'b11111110111101010000001111100110;
   assign mem[270687:270656] = 32'b11111111010011101011110011010011;
   assign mem[270719:270688] = 32'b11111001000000001100000111000000;
   assign mem[270751:270720] = 32'b11111001101001111011010110101000;
   assign mem[270783:270752] = 32'b11110111000010110111101000110000;
   assign mem[270815:270784] = 32'b11111011111100111010001010010000;
   assign mem[270847:270816] = 32'b00000100001111111011110110110000;
   assign mem[270879:270848] = 32'b00000010010001101001110000001000;
   assign mem[270911:270880] = 32'b11111011110011010110110011111000;
   assign mem[270943:270912] = 32'b00000010010010101001101101000100;
   assign mem[270975:270944] = 32'b11111110001011010111000000010100;
   assign mem[271007:270976] = 32'b00000010000001101000111011111000;
   assign mem[271039:271008] = 32'b00000011110010100011011111010000;
   assign mem[271071:271040] = 32'b00000010111111111000011000101100;
   assign mem[271103:271072] = 32'b11111101111110101111100110011100;
   assign mem[271135:271104] = 32'b00000101011110000011100110000000;
   assign mem[271167:271136] = 32'b11111101110011110010010110001100;
   assign mem[271199:271168] = 32'b00000010111110110000101101000100;
   assign mem[271231:271200] = 32'b11110110111101000101001110000000;
   assign mem[271263:271232] = 32'b11111001001111100111111100001000;
   assign mem[271295:271264] = 32'b00000011110010000000111101001000;
   assign mem[271327:271296] = 32'b00000000010010011111110011110010;
   assign mem[271359:271328] = 32'b11111010000011100100111101010000;
   assign mem[271391:271360] = 32'b11110011111110101000110101000000;
   assign mem[271423:271392] = 32'b11110111110111100101110010010000;
   assign mem[271455:271424] = 32'b11111101011001111011111000011100;
   assign mem[271487:271456] = 32'b00000110100011001101011000010000;
   assign mem[271519:271488] = 32'b00001011100101011110010000000000;
   assign mem[271551:271520] = 32'b11110111111001011100100000100000;
   assign mem[271583:271552] = 32'b11110101111111000010110011100000;
   assign mem[271615:271584] = 32'b11111111010001111010111110000011;
   assign mem[271647:271616] = 32'b00001000010010010110101011110000;
   assign mem[271679:271648] = 32'b00000111100110111011001010111000;
   assign mem[271711:271680] = 32'b11110110111011101010111001110000;
   assign mem[271743:271712] = 32'b11111011100110100110100110100000;
   assign mem[271775:271744] = 32'b11111101110001110110000111011100;
   assign mem[271807:271776] = 32'b00000010001101000111100010001100;
   assign mem[271839:271808] = 32'b00000111110101011111011111111000;
   assign mem[271871:271840] = 32'b00000000100111101010111011101011;
   assign mem[271903:271872] = 32'b11111111000110111010011110011101;
   assign mem[271935:271904] = 32'b11111100110111100100100011001000;
   assign mem[271967:271936] = 32'b11111101001000101110000101111100;
   assign mem[271999:271968] = 32'b00000100101110001110001111100000;
   assign mem[272031:272000] = 32'b11111101001001001110010011010100;
   assign mem[272063:272032] = 32'b11110110011100110001011101010000;
   assign mem[272095:272064] = 32'b11111001101110001000100001010000;
   assign mem[272127:272096] = 32'b00000100011010001011111010001000;
   assign mem[272159:272128] = 32'b11110001000000101101010100010000;
   assign mem[272191:272160] = 32'b00000111100101000011010000011000;
   assign mem[272223:272192] = 32'b00001000010011111010000001000000;
   assign mem[272255:272224] = 32'b11111011110100100100110000001000;
   assign mem[272287:272256] = 32'b11111111000000110110010111011000;
   assign mem[272319:272288] = 32'b00000000011001001001000011000101;
   assign mem[272351:272320] = 32'b11111110110110000101010011011000;
   assign mem[272383:272352] = 32'b11101000100110100010100111100000;
   assign mem[272415:272384] = 32'b11111100101000001000001110010000;
   assign mem[272447:272416] = 32'b00000110100011101101111001101000;
   assign mem[272479:272448] = 32'b11111010101101001001011111010000;
   assign mem[272511:272480] = 32'b11111011110010100100011110110000;
   assign mem[272543:272512] = 32'b00000110101010101100010100110000;
   assign mem[272575:272544] = 32'b11111111110001100011001010000111;
   assign mem[272607:272576] = 32'b00000000000010000001011011110011;
   assign mem[272639:272608] = 32'b00000010010000011110001001101000;
   assign mem[272671:272640] = 32'b00000010001001010101010000011100;
   assign mem[272703:272672] = 32'b00000001111100111000110000010010;
   assign mem[272735:272704] = 32'b00000100010000011100111011110000;
   assign mem[272767:272736] = 32'b11110101011100011010100001100000;
   assign mem[272799:272768] = 32'b00000010101010101101010011011100;
   assign mem[272831:272800] = 32'b11111101110000110011100101001100;
   assign mem[272863:272832] = 32'b11111011011011000010101100110000;
   assign mem[272895:272864] = 32'b00000101011000110010110010111000;
   assign mem[272927:272896] = 32'b11110110001011011110101100000000;
   assign mem[272959:272928] = 32'b00000000010000000010011100001101;
   assign mem[272991:272960] = 32'b11111000000110101011001001111000;
   assign mem[273023:272992] = 32'b11111010001011101001011000011000;
   assign mem[273055:273024] = 32'b11111101110110100111010000101000;
   assign mem[273087:273056] = 32'b00000010000101001000000001101000;
   assign mem[273119:273088] = 32'b11111010001001100100111000010000;
   assign mem[273151:273120] = 32'b00000001000010010010011100111110;
   assign mem[273183:273152] = 32'b00000100101010111110001111100000;
   assign mem[273215:273184] = 32'b11111110110100000110111011110100;
   assign mem[273247:273216] = 32'b00000111001100000010111010100000;
   assign mem[273279:273248] = 32'b00000110010101000011110000100000;
   assign mem[273311:273280] = 32'b11111100001110010010100101101000;
   assign mem[273343:273312] = 32'b11111110101011111100010011011100;
   assign mem[273375:273344] = 32'b00000010011001101101101000101100;
   assign mem[273407:273376] = 32'b00001001011010110011110100110000;
   assign mem[273439:273408] = 32'b11111101101100001101001010111100;
   assign mem[273471:273440] = 32'b11110000010000010000110100100000;
   assign mem[273503:273472] = 32'b11111001100110010001110111000000;
   assign mem[273535:273504] = 32'b00000010011011100100111011000000;
   assign mem[273567:273536] = 32'b00000101010110110111010000010000;
   assign mem[273599:273568] = 32'b00000001010011100101110011001010;
   assign mem[273631:273600] = 32'b00000100111101101100100001101000;
   assign mem[273663:273632] = 32'b00000000100101110111011100111111;
   assign mem[273695:273664] = 32'b11111100010011011111011111111100;
   assign mem[273727:273696] = 32'b00000001001010101110011100010110;
   assign mem[273759:273728] = 32'b00001001000011100111100000100000;
   assign mem[273791:273760] = 32'b00000000000000111011100100101010;
   assign mem[273823:273792] = 32'b11110111011010111110000100100000;
   assign mem[273855:273824] = 32'b00000101110001110100101010001000;
   assign mem[273887:273856] = 32'b11111111010010100000001111111000;
   assign mem[273919:273888] = 32'b00000000100110110100100101110110;
   assign mem[273951:273920] = 32'b00001010010011100110100000000000;
   assign mem[273983:273952] = 32'b11111111110110011100100010101011;
   assign mem[274015:273984] = 32'b00000010011000011001110100000100;
   assign mem[274047:274016] = 32'b11111110001110111001010111110010;
   assign mem[274079:274048] = 32'b00000011011011110000000111100000;
   assign mem[274111:274080] = 32'b11111110111101101111101011110110;
   assign mem[274143:274112] = 32'b11111100010011100000011110001100;
   assign mem[274175:274144] = 32'b00000101110000010010011111110000;
   assign mem[274207:274176] = 32'b11111011111011110001010111001000;
   assign mem[274239:274208] = 32'b00000000000111001111110110001010;
   assign mem[274271:274240] = 32'b11111000010111100000000100000000;
   assign mem[274303:274272] = 32'b00000000001010011111011100010011;
   assign mem[274335:274304] = 32'b00000001000110100101011011000010;
   assign mem[274367:274336] = 32'b00000001011110010111101101010000;
   assign mem[274399:274368] = 32'b11111100110010111101001101110100;
   assign mem[274431:274400] = 32'b11111110000110100010011100101100;
   assign mem[274463:274432] = 32'b11111001100001111100010011111000;
   assign mem[274495:274464] = 32'b00000010111111100011000101100000;
   assign mem[274527:274496] = 32'b11111111000100101110011100100110;
   assign mem[274559:274528] = 32'b00000011100010000001100111011000;
   assign mem[274591:274560] = 32'b00000010000110110011001001000000;
   assign mem[274623:274592] = 32'b00000010111110101000000001110100;
   assign mem[274655:274624] = 32'b11111101111100000010001100001100;
   assign mem[274687:274656] = 32'b11111011000011010101111001011000;
   assign mem[274719:274688] = 32'b00000100101010101010000110010000;
   assign mem[274751:274720] = 32'b11110101000111111010001011000000;
   assign mem[274783:274752] = 32'b11111011111011011000101110011000;
   assign mem[274815:274784] = 32'b00000001101111000101010111010000;
   assign mem[274847:274816] = 32'b00000000011010001011010110100110;
   assign mem[274879:274848] = 32'b11111110101000011011001011100110;
   assign mem[274911:274880] = 32'b11111110100011011011111110110100;
   assign mem[274943:274912] = 32'b11111111011001000111000101110110;
   assign mem[274975:274944] = 32'b00001001000000011011000000000000;
   assign mem[275007:274976] = 32'b11101100011101100001101010100000;
   assign mem[275039:275008] = 32'b00000011001000001100111000100000;
   assign mem[275071:275040] = 32'b11111110110000100001000111110010;
   assign mem[275103:275072] = 32'b00000010000111010001100001111100;
   assign mem[275135:275104] = 32'b11111001111001001000101101010000;
   assign mem[275167:275136] = 32'b00000111111011000000101101110000;
   assign mem[275199:275168] = 32'b11111100101011000011011010001100;
   assign mem[275231:275200] = 32'b11110100010010101110001001000000;
   assign mem[275263:275232] = 32'b11101101001010100001100010100000;
   assign mem[275295:275264] = 32'b11111100010100110011110110000000;
   assign mem[275327:275296] = 32'b00000100000100011101000110000000;
   assign mem[275359:275328] = 32'b00000110000111100100101100110000;
   assign mem[275391:275360] = 32'b11110110101001000011001010110000;
   assign mem[275423:275392] = 32'b00000010111001000000000000001000;
   assign mem[275455:275424] = 32'b11111100110101001110000010001100;
   assign mem[275487:275456] = 32'b00000100011111101100010100001000;
   assign mem[275519:275488] = 32'b00000011110000010111010100011100;
   assign mem[275551:275520] = 32'b11110110100001010111100111000000;
   assign mem[275583:275552] = 32'b11111010001101000100111101101000;
   assign mem[275615:275584] = 32'b00001001010011101111001000110000;
   assign mem[275647:275616] = 32'b11111100110101000100011011100000;
   assign mem[275679:275648] = 32'b11110110010010011110011010100000;
   assign mem[275711:275680] = 32'b00000110100111010111000000110000;
   assign mem[275743:275712] = 32'b00001110110001011110111101100000;
   assign mem[275775:275744] = 32'b11111111011100010001110010001000;
   assign mem[275807:275776] = 32'b11110101110110111000101001000000;
   assign mem[275839:275808] = 32'b11111011101011110000000110101000;
   assign mem[275871:275840] = 32'b00000101100011001111000100110000;
   assign mem[275903:275872] = 32'b00000110011100001001100111001000;
   assign mem[275935:275904] = 32'b00000000011010011011001010111000;
   assign mem[275967:275936] = 32'b11111101100001110100000100110100;
   assign mem[275999:275968] = 32'b00000000111111011010011000000010;
   assign mem[276031:276000] = 32'b11111111110111010110010110011011;
   assign mem[276063:276032] = 32'b11110001011110110000101110010000;
   assign mem[276095:276064] = 32'b00000100010110100000011010101000;
   assign mem[276127:276096] = 32'b11111110010010101011101100000010;
   assign mem[276159:276128] = 32'b11111110010001110010110100110100;
   assign mem[276191:276160] = 32'b00000011001010101011101010111100;
   assign mem[276223:276192] = 32'b11101110000110110011010000100000;
   assign mem[276255:276224] = 32'b11110110110010001100010001100000;
   assign mem[276287:276256] = 32'b00000010111010011001101010111100;
   assign mem[276319:276288] = 32'b00000001001111110000101100011110;
   assign mem[276351:276320] = 32'b11111110000011011101111101001010;
   assign mem[276383:276352] = 32'b00000000101000010000001110101010;
   assign mem[276415:276384] = 32'b00001011100110010011100110100000;
   assign mem[276447:276416] = 32'b00000100001011101000110100010000;
   assign mem[276479:276448] = 32'b11111010011110100111000010111000;
   assign mem[276511:276480] = 32'b11110010001010101010010000110000;
   assign mem[276543:276512] = 32'b00000111111010010010110000011000;
   assign mem[276575:276544] = 32'b00000000100010001100100110001011;
   assign mem[276607:276576] = 32'b00001010100010000010001110000000;
   assign mem[276639:276608] = 32'b11111111011110100101100010101110;
   assign mem[276671:276640] = 32'b11101000010011000001010101000000;
   assign mem[276703:276672] = 32'b11111011000111101010111011011000;
   assign mem[276735:276704] = 32'b11111110100100110111101111010100;
   assign mem[276767:276736] = 32'b00000101001010101001001111011000;
   assign mem[276799:276768] = 32'b00000010001100010110001001001100;
   assign mem[276831:276800] = 32'b11111101111111011011110101110000;
   assign mem[276863:276832] = 32'b00000011101000001101010000101100;
   assign mem[276895:276864] = 32'b00000100111111001000111111001000;
   assign mem[276927:276896] = 32'b11110101001100001100100010110000;
   assign mem[276959:276928] = 32'b11111111010000001101100101001100;
   assign mem[276991:276960] = 32'b11111000111000010100000001101000;
   assign mem[277023:276992] = 32'b11111110110010100111010001100100;
   assign mem[277055:277024] = 32'b00000111100100101111001000111000;
   assign mem[277087:277056] = 32'b00000101000000110010000111000000;
   assign mem[277119:277088] = 32'b11110111110000011110000101010000;
   assign mem[277151:277120] = 32'b11110110110001001100000100110000;
   assign mem[277183:277152] = 32'b11111110110011000000110001000010;
   assign mem[277215:277184] = 32'b11111100000110001001110111101100;
   assign mem[277247:277216] = 32'b00000101100111111111010110110000;
   assign mem[277279:277248] = 32'b00000010001110001111011011001100;
   assign mem[277311:277280] = 32'b00000001110110110111110100010100;
   assign mem[277343:277312] = 32'b11111111111100010011000100101001;
   assign mem[277375:277344] = 32'b00000110001111010111010001001000;
   assign mem[277407:277376] = 32'b11111111111010001101000001100000;
   assign mem[277439:277408] = 32'b11111001011010011110111111100000;
   assign mem[277471:277440] = 32'b00000101010001001100011000110000;
   assign mem[277503:277472] = 32'b00000101010100101010110111111000;
   assign mem[277535:277504] = 32'b00000100001111011011001111111000;
   assign mem[277567:277536] = 32'b11111001001101100001100010001000;
   assign mem[277599:277568] = 32'b11111001010000000000100001110000;
   assign mem[277631:277600] = 32'b11110101111101100011010001000000;
   assign mem[277663:277632] = 32'b11111100111001110111100011010100;
   assign mem[277695:277664] = 32'b00000000010110110110100101010000;
   assign mem[277727:277696] = 32'b11111100000011011110000000001000;
   assign mem[277759:277728] = 32'b00000011111011010100000100001000;
   assign mem[277791:277760] = 32'b11110111111110001011100100100000;
   assign mem[277823:277792] = 32'b11101110001110111100000010100000;
   assign mem[277855:277824] = 32'b00000100000100010000001100001000;
   assign mem[277887:277856] = 32'b00000111000001100100011011111000;
   assign mem[277919:277888] = 32'b11111101111010000110111110011000;
   assign mem[277951:277920] = 32'b00000110010010000010010011000000;
   assign mem[277983:277952] = 32'b00001010011001000110010001000000;
   assign mem[278015:277984] = 32'b11101111011001110100111101100000;
   assign mem[278047:278016] = 32'b00000001010001111010000101010000;
   assign mem[278079:278048] = 32'b11110111000110000110001100100000;
   assign mem[278111:278080] = 32'b11111000001011000111111010110000;
   assign mem[278143:278112] = 32'b11111011110110000010111111011000;
   assign mem[278175:278144] = 32'b11111001001001000110010100010000;
   assign mem[278207:278176] = 32'b00000001111011111110001011100000;
   assign mem[278239:278208] = 32'b11111100011011111110111011111000;
   assign mem[278271:278240] = 32'b00000100100001101110110000001000;
   assign mem[278303:278272] = 32'b00000110111010100110101000111000;
   assign mem[278335:278304] = 32'b11111010100000110101100011001000;
   assign mem[278367:278336] = 32'b00000001010010101110110000010000;
   assign mem[278399:278368] = 32'b11111111010001110010111101111101;
   assign mem[278431:278400] = 32'b11111101100010001100101110000000;
   assign mem[278463:278432] = 32'b11111110110101000110010100110110;
   assign mem[278495:278464] = 32'b11111011101010000110100001110000;
   assign mem[278527:278496] = 32'b00000101000100001010000001111000;
   assign mem[278559:278528] = 32'b00000100010111010010000010000000;
   assign mem[278591:278560] = 32'b11110101011000001110010110000000;
   assign mem[278623:278592] = 32'b11110101011101100001010010100000;
   assign mem[278655:278624] = 32'b00001001100010110001000000000000;
   assign mem[278687:278656] = 32'b00001001101011001000011011110000;
   assign mem[278719:278688] = 32'b00000100100100001000100111111000;
   assign mem[278751:278720] = 32'b11111001111110010110010000111000;
   assign mem[278783:278752] = 32'b11110111101111010111010000000000;
   assign mem[278815:278784] = 32'b00000011100000101111111011001100;
   assign mem[278847:278816] = 32'b11111110111010010011011011011010;
   assign mem[278879:278848] = 32'b11110110011101100100010001000000;
   assign mem[278911:278880] = 32'b11111100111111010101111100100000;
   assign mem[278943:278912] = 32'b11111110010001110111111000101000;
   assign mem[278975:278944] = 32'b11111110100000101111101011010110;
   assign mem[279007:278976] = 32'b00000111110000110011011010110000;
   assign mem[279039:279008] = 32'b00000010100010101000111100101100;
   assign mem[279071:279040] = 32'b00000000110000001100011101100001;
   assign mem[279103:279072] = 32'b00000100011101101010000011000000;
   assign mem[279135:279104] = 32'b11110111110000000101100111100000;
   assign mem[279167:279136] = 32'b00000010101100011111101101101100;
   assign mem[279199:279168] = 32'b11111111101011100011101111010011;
   assign mem[279231:279200] = 32'b00000100011111011100001011010000;
   assign mem[279263:279232] = 32'b11111101111100000111001100011100;
   assign mem[279295:279264] = 32'b00000011110101011111011100010100;
   assign mem[279327:279296] = 32'b11111111011001100000011001011100;
   assign mem[279359:279328] = 32'b11111111111000100001000011011110;
   assign mem[279391:279360] = 32'b11111100010111101111001010010100;
   assign mem[279423:279392] = 32'b11111010111001010011001100100000;
   assign mem[279455:279424] = 32'b11111001111000011110100000000000;
   assign mem[279487:279456] = 32'b00000111010010111110000000001000;
   assign mem[279519:279488] = 32'b00000001110011000011111010010110;
   assign mem[279551:279520] = 32'b11111111100110011110110010000101;
   assign mem[279583:279552] = 32'b11110111100011000110100110100000;
   assign mem[279615:279584] = 32'b11111011110101110101111000010000;
   assign mem[279647:279616] = 32'b00000100000111011101101100100000;
   assign mem[279679:279648] = 32'b00001010110111010011001111000000;
   assign mem[279711:279680] = 32'b00001100100110011110100010100000;
   assign mem[279743:279712] = 32'b11111111110000000001001110110100;
   assign mem[279775:279744] = 32'b11101101100011101111100100100000;
   assign mem[279807:279776] = 32'b11111110110001110101100011100010;
   assign mem[279839:279808] = 32'b11101111101110011010101100100000;
   assign mem[279871:279840] = 32'b00000110100010000100010100000000;
   assign mem[279903:279872] = 32'b11111010011110111010110001111000;
   assign mem[279935:279904] = 32'b00010000011001100000111000000000;
   assign mem[279967:279936] = 32'b11110001000110011001101011100000;
   assign mem[279999:279968] = 32'b11111101111010000001100011001000;
   assign mem[280031:280000] = 32'b00000001011110110100000001011000;
   assign mem[280063:280032] = 32'b00000010100000001010111110000100;
   assign mem[280095:280064] = 32'b00000000100101010111011110010111;
   assign mem[280127:280096] = 32'b11111111000000000000001111011011;
   assign mem[280159:280128] = 32'b11111110101011010010101010100100;
   assign mem[280191:280160] = 32'b11111000011111000000100001101000;
   assign mem[280223:280192] = 32'b11111100011100101111001111011000;
   assign mem[280255:280224] = 32'b11111110100011111100110011001110;
   assign mem[280287:280256] = 32'b11111100011101000010010110100000;
   assign mem[280319:280288] = 32'b00000001111010101001111001010000;
   assign mem[280351:280320] = 32'b11111001000000010100010010100000;
   assign mem[280383:280352] = 32'b00000101101110010101101101010000;
   assign mem[280415:280384] = 32'b11111011111001001111000101000000;
   assign mem[280447:280416] = 32'b00000010011010011100010101000100;
   assign mem[280479:280448] = 32'b00001010100101101111001000110000;
   assign mem[280511:280480] = 32'b11111001000000000000101110011000;
   assign mem[280543:280512] = 32'b11110110000110100000001010100000;
   assign mem[280575:280544] = 32'b00001010000100011100010000110000;
   assign mem[280607:280576] = 32'b11111000000100010001000110001000;
   assign mem[280639:280608] = 32'b11111110101100011000101010011010;
   assign mem[280671:280640] = 32'b00000000001000101001000001011011;
   assign mem[280703:280672] = 32'b11111110111101111011011110001010;
   assign mem[280735:280704] = 32'b00000010011100110111101100101000;
   assign mem[280767:280736] = 32'b00000100010110111110011111011000;
   assign mem[280799:280768] = 32'b11111011000111000000011001010000;
   assign mem[280831:280800] = 32'b00000100100000110010000110001000;
   assign mem[280863:280832] = 32'b00000110010111011100001111111000;
   assign mem[280895:280864] = 32'b11111000000001101111001110011000;
   assign mem[280927:280896] = 32'b00000000101111000101000110000011;
   assign mem[280959:280928] = 32'b11111111101101000111110111010110;
   assign mem[280991:280960] = 32'b11111111110100000100010100001111;
   assign mem[281023:280992] = 32'b11111011010111011000110100111000;
   assign mem[281055:281024] = 32'b00000001001000000011001010001000;
   assign mem[281087:281056] = 32'b11111110101001011100101011010100;
   assign mem[281119:281088] = 32'b11111111111101001011111110001010;
   assign mem[281151:281120] = 32'b00000010100100111100001100110000;
   assign mem[281183:281152] = 32'b11110111101111110000011100110000;
   assign mem[281215:281184] = 32'b00001000001001011000000110000000;
   assign mem[281247:281216] = 32'b11111001010101000010111010101000;
   assign mem[281279:281248] = 32'b11111001111101010100100000010000;
   assign mem[281311:281280] = 32'b00000100001011110001000101110000;
   assign mem[281343:281312] = 32'b00000000000110110010111111000000;
   assign mem[281375:281344] = 32'b00000000111101011101100100100000;
   assign mem[281407:281376] = 32'b11111100001111100100000001110000;
   assign mem[281439:281408] = 32'b00000010010011110010011100111100;
   assign mem[281471:281440] = 32'b00000010101100111101011011110100;
   assign mem[281503:281472] = 32'b00000010100111101111010111111100;
   assign mem[281535:281504] = 32'b11111101100011101010111010010100;
   assign mem[281567:281536] = 32'b00000001111101100110110110110100;
   assign mem[281599:281568] = 32'b11111100011111010100110011010100;
   assign mem[281631:281600] = 32'b11110110111001001010101100010000;
   assign mem[281663:281632] = 32'b00000111000011000001111000101000;
   assign mem[281695:281664] = 32'b11111110001011110011000001111110;
   assign mem[281727:281696] = 32'b00000111000111101001010001101000;
   assign mem[281759:281728] = 32'b00000010100101110000000001100000;
   assign mem[281791:281760] = 32'b11111101101010110111110000100000;
   assign mem[281823:281792] = 32'b00000000111100000010010100001001;
   assign mem[281855:281824] = 32'b00000000111110001101100011001100;
   assign mem[281887:281856] = 32'b00000001000100010011110000010110;
   assign mem[281919:281888] = 32'b00001001001010101111111001100000;
   assign mem[281951:281920] = 32'b11111111111000101010010100011111;
   assign mem[281983:281952] = 32'b00000000101011111011110101110100;
   assign mem[282015:281984] = 32'b11111101101110111011111000011000;
   assign mem[282047:282016] = 32'b11110100110110110110000011100000;
   assign mem[282079:282048] = 32'b00000000110110001000000111001010;
   assign mem[282111:282080] = 32'b11110100011000110110110010110000;
   assign mem[282143:282112] = 32'b00000011010010111000100111011000;
   assign mem[282175:282144] = 32'b11111111101111011000111001101011;
   assign mem[282207:282176] = 32'b00000101100100111110010001100000;
   assign mem[282239:282208] = 32'b00000010000100100101100111000100;
   assign mem[282271:282240] = 32'b11111111011010111100011111011010;
   assign mem[282303:282272] = 32'b11111011010110010110001010011000;
   assign mem[282335:282304] = 32'b00000000100000111011001001001101;
   assign mem[282367:282336] = 32'b00000000110011011001010111101110;
   assign mem[282399:282368] = 32'b00000001000100001101111111010110;
   assign mem[282431:282400] = 32'b11110000100100001100000001100000;
   assign mem[282463:282432] = 32'b11111011000001011011011011101000;
   assign mem[282495:282464] = 32'b00000010010011001001111010011100;
   assign mem[282527:282496] = 32'b00000100100111001000100011100000;
   assign mem[282559:282528] = 32'b00000000101011011000100111101101;
   assign mem[282591:282560] = 32'b00000000001111101111100001100001;
   assign mem[282623:282592] = 32'b00000111100101111100010001001000;
   assign mem[282655:282624] = 32'b00010000100001100110100001100000;
   assign mem[282687:282656] = 32'b11101111001100110111111110000000;
   assign mem[282719:282688] = 32'b00001111100111011001100001010000;
   assign mem[282751:282720] = 32'b00000011111001100011101100110100;
   assign mem[282783:282752] = 32'b11101111000010100010110100000000;
   assign mem[282815:282784] = 32'b00000010110111010001011001001000;
   assign mem[282847:282816] = 32'b11110011010100000000111101010000;
   assign mem[282879:282848] = 32'b11111011101001100111010000010000;
   assign mem[282911:282880] = 32'b11110110001101110011011000010000;
   assign mem[282943:282912] = 32'b11110101001001101000111111010000;
   assign mem[282975:282944] = 32'b11111100110011001011111100110100;
   assign mem[283007:282976] = 32'b00000111100111000000100101011000;
   assign mem[283039:283008] = 32'b11111111001101011010000011011011;
   assign mem[283071:283040] = 32'b00000000111001011010001001110000;
   assign mem[283103:283072] = 32'b00000101100111011000110000101000;
   assign mem[283135:283104] = 32'b00000100001010011010100000100000;
   assign mem[283167:283136] = 32'b11111100010011101111110010101000;
   assign mem[283199:283168] = 32'b00000010110101011001101001101100;
   assign mem[283231:283200] = 32'b11110010011110010101010001010000;
   assign mem[283263:283232] = 32'b11110011011110110001000101000000;
   assign mem[283295:283264] = 32'b00000000011110000001111110010011;
   assign mem[283327:283296] = 32'b00000101100101001000000001111000;
   assign mem[283359:283328] = 32'b11111100100101010010010001100000;
   assign mem[283391:283360] = 32'b00000010100101101100111010100000;
   assign mem[283423:283392] = 32'b00000101011000100010011110101000;
   assign mem[283455:283424] = 32'b11111101001110100011101011101100;
   assign mem[283487:283456] = 32'b11111111010001000010111011010001;
   assign mem[283519:283488] = 32'b00000001101001111001101110010010;
   assign mem[283551:283520] = 32'b11101110001000100111010010100000;
   assign mem[283583:283552] = 32'b00000001100100000000111001100110;
   assign mem[283615:283584] = 32'b11111111011011000011111100010011;
   assign mem[283647:283616] = 32'b00000011111111011111110001100100;
   assign mem[283679:283648] = 32'b00000001000001010011110010100110;
   assign mem[283711:283680] = 32'b11111001110100100010000110010000;
   assign mem[283743:283712] = 32'b11110111111111111001100100010000;
   assign mem[283775:283744] = 32'b11111100000111011001111111111100;
   assign mem[283807:283776] = 32'b00000011010110011000100001000000;
   assign mem[283839:283808] = 32'b00000011000010000100101110000000;
   assign mem[283871:283840] = 32'b11111110110000010100110001010110;
   assign mem[283903:283872] = 32'b00000001000011110011111011011010;
   assign mem[283935:283904] = 32'b00000100000010000000101010111000;
   assign mem[283967:283936] = 32'b00000010110010001011110011101100;
   assign mem[283999:283968] = 32'b11111010111111001101000100111000;
   assign mem[284031:284000] = 32'b11111010000011011101100011110000;
   assign mem[284063:284032] = 32'b11111101011110010010011100010000;
   assign mem[284095:284064] = 32'b00000001010010011011010111100110;
   assign mem[284127:284096] = 32'b11111110000111001111000010011010;
   assign mem[284159:284128] = 32'b11111111110100100111110001010000;
   assign mem[284191:284160] = 32'b11111011101000010110111101010000;
   assign mem[284223:284192] = 32'b00000011110010101010110000011100;
   assign mem[284255:284224] = 32'b11111110010001001010101110101000;
   assign mem[284287:284256] = 32'b00000000100000111001101110110010;
   assign mem[284319:284288] = 32'b00000010111000010101111010110100;
   assign mem[284351:284320] = 32'b00000001010000010111100011100000;
   assign mem[284383:284352] = 32'b11111011011000100010110011000000;
   assign mem[284415:284384] = 32'b11111011000000101011001101110000;
   assign mem[284447:284416] = 32'b11110010101101110110111100000000;
   assign mem[284479:284448] = 32'b00001001111011110101110111110000;
   assign mem[284511:284480] = 32'b00000111110100101010110110001000;
   assign mem[284543:284512] = 32'b11110011110010001110000100100000;
   assign mem[284575:284544] = 32'b11111001010001011010010011000000;
   assign mem[284607:284576] = 32'b00000011000101101101010010001100;
   assign mem[284639:284608] = 32'b11110110101101011010010100010000;
   assign mem[284671:284640] = 32'b00000010001101100111010100000100;
   assign mem[284703:284672] = 32'b11111111000011101111101111110101;
   assign mem[284735:284704] = 32'b00000101001000010011011000111000;
   assign mem[284767:284736] = 32'b00000011011010100101011000010000;
   assign mem[284799:284768] = 32'b11111110100100010011010110101110;
   assign mem[284831:284800] = 32'b11111010011011011010011100010000;
   assign mem[284863:284832] = 32'b00000111110100100110011001010000;
   assign mem[284895:284864] = 32'b00000100001111000111010110111000;
   assign mem[284927:284896] = 32'b11111000001001000100001000100000;
   assign mem[284959:284928] = 32'b00000000111101010010100101001111;
   assign mem[284991:284960] = 32'b00000001101001101111010111110110;
   assign mem[285023:284992] = 32'b00001000000110010010010101100000;
   assign mem[285055:285024] = 32'b11111000001111010101001010010000;
   assign mem[285087:285056] = 32'b11110001001100011110010111000000;
   assign mem[285119:285088] = 32'b11111110101011000001011001111110;
   assign mem[285151:285120] = 32'b11111011010001000111010100111000;
   assign mem[285183:285152] = 32'b11111011011100001110101110010000;
   assign mem[285215:285184] = 32'b11111100010010000100000110111100;
   assign mem[285247:285216] = 32'b11111110000001001100011100001010;
   assign mem[285279:285248] = 32'b00000010011010011000111011110000;
   assign mem[285311:285280] = 32'b00000010111000100110110001001100;
   assign mem[285343:285312] = 32'b00000101010101011111000110011000;
   assign mem[285375:285344] = 32'b11111100010111000110110010001100;
   assign mem[285407:285376] = 32'b00000011111110010010101001000000;
   assign mem[285439:285408] = 32'b00000000001101010011111110001111;
   assign mem[285471:285440] = 32'b11111110000110000110001011100010;
   assign mem[285503:285472] = 32'b11111010110100100001010111000000;
   assign mem[285535:285504] = 32'b00000000001110110010100011010011;
   assign mem[285567:285536] = 32'b00000000001000001010110001101100;
   assign mem[285599:285568] = 32'b11111010100011100100010110110000;
   assign mem[285631:285600] = 32'b11111011101010110110110101000000;
   assign mem[285663:285632] = 32'b00000100000010111011000110001000;
   assign mem[285695:285664] = 32'b11110111111000111010110010010000;
   assign mem[285727:285696] = 32'b00000110101011001100011100101000;
   assign mem[285759:285728] = 32'b00000011001011000110001101001100;
   assign mem[285791:285760] = 32'b11110110011110000001100101010000;
   assign mem[285823:285792] = 32'b00000101011100110110011000100000;
   assign mem[285855:285824] = 32'b00000011011010011111001101011100;
   assign mem[285887:285856] = 32'b11110011111000110011000101000000;
   assign mem[285919:285888] = 32'b00000101001111010000101100010000;
   assign mem[285951:285920] = 32'b11110111111011101101111100010000;
   assign mem[285983:285952] = 32'b00000101100011011001111100110000;
   assign mem[286015:285984] = 32'b00000100100011011111011010000000;
   assign mem[286047:286016] = 32'b00000110111010110101011000000000;
   assign mem[286079:286048] = 32'b11111100100111101111100101000000;
   assign mem[286111:286080] = 32'b00000111101111001101101100101000;
   assign mem[286143:286112] = 32'b00000000111011010111010000100000;
   assign mem[286175:286144] = 32'b00000101001011111010110010101000;
   assign mem[286207:286176] = 32'b11101010011011100101100110100000;
   assign mem[286239:286208] = 32'b00001011000000000010010000010000;
   assign mem[286271:286240] = 32'b11111100001000001000110000101000;
   assign mem[286303:286272] = 32'b11110111110110001111111010110000;
   assign mem[286335:286304] = 32'b00000110011000111000011110000000;
   assign mem[286367:286336] = 32'b11100110001001001100110001100000;
   assign mem[286399:286368] = 32'b11111110000001110101100010011010;
   assign mem[286431:286400] = 32'b00000000011001001101101000101110;
   assign mem[286463:286432] = 32'b00000001101101101001001101111100;
   assign mem[286495:286464] = 32'b00000110000111100111001001011000;
   assign mem[286527:286496] = 32'b11110100000100110011011011100000;
   assign mem[286559:286528] = 32'b00001010101111011010010101110000;
   assign mem[286591:286560] = 32'b11111110010100000011000101111000;
   assign mem[286623:286592] = 32'b11110010100010010011111011110000;
   assign mem[286655:286624] = 32'b00000011010111001101101010000100;
   assign mem[286687:286656] = 32'b11111011010001011010101100101000;
   assign mem[286719:286688] = 32'b11111111011100011110011111100111;
   assign mem[286751:286720] = 32'b11111111111000011111100111100010;
   assign mem[286783:286752] = 32'b11111000010110011010100010100000;
   assign mem[286815:286784] = 32'b00000110010111001001011100010000;
   assign mem[286847:286816] = 32'b00001100011111010111010110000000;
   assign mem[286879:286848] = 32'b00000000001010000010101111000111;
   assign mem[286911:286880] = 32'b11111001010001110011100010101000;
   assign mem[286943:286912] = 32'b00000011011111011000000010000100;
   assign mem[286975:286944] = 32'b11111101101001100011011110001100;
   assign mem[287007:286976] = 32'b00000111110001101101001111111000;
   assign mem[287039:287008] = 32'b11101001011110100000000010000000;
   assign mem[287071:287040] = 32'b11111011101010000100001011110000;
   assign mem[287103:287072] = 32'b11111100000000111000001010110000;
   assign mem[287135:287104] = 32'b11111011001111000111111111010000;
   assign mem[287167:287136] = 32'b00000001010101011000011110101100;
   assign mem[287199:287168] = 32'b11111110001000101111110111100110;
   assign mem[287231:287200] = 32'b00000100000000010010111011100000;
   assign mem[287263:287232] = 32'b00000011010010111001000110100100;
   assign mem[287295:287264] = 32'b11111100101001001010111111000100;
   assign mem[287327:287296] = 32'b11111011000110001011001001001000;
   assign mem[287359:287328] = 32'b00000000011000000000111111111101;
   assign mem[287391:287360] = 32'b00000001111111101100100111010010;
   assign mem[287423:287392] = 32'b11111010000111100011101010110000;
   assign mem[287455:287424] = 32'b11110101001010000100000101000000;
   assign mem[287487:287456] = 32'b00000010001001010011000001010000;
   assign mem[287519:287488] = 32'b11111000110011100101111101011000;
   assign mem[287551:287520] = 32'b00000100100011000000010010011000;
   assign mem[287583:287552] = 32'b00000011001001011000000000110100;
   assign mem[287615:287584] = 32'b11111111010001100111100100011010;
   assign mem[287647:287616] = 32'b00000010100111010011000110100000;
   assign mem[287679:287648] = 32'b11110010111001101111011111000000;
   assign mem[287711:287680] = 32'b00000011001101001001011000100000;
   assign mem[287743:287712] = 32'b00000000100110110000101110001100;
   assign mem[287775:287744] = 32'b11111011010000100110010110101000;
   assign mem[287807:287776] = 32'b00000001001110111110011110100000;
   assign mem[287839:287808] = 32'b00000001110011010000111100110010;
   assign mem[287871:287840] = 32'b00001011100010110100111011010000;
   assign mem[287903:287872] = 32'b11111000000001000010101101100000;
   assign mem[287935:287904] = 32'b11111001010000010110001110101000;
   assign mem[287967:287936] = 32'b11111101100110100001101000100100;
   assign mem[287999:287968] = 32'b11111010001110111011111111011000;
   assign mem[288031:288000] = 32'b11101011110011101100110010000000;
   assign mem[288063:288032] = 32'b00000011001101011011011011110100;
   assign mem[288095:288064] = 32'b11111101101011010111101101110000;
   assign mem[288127:288096] = 32'b11111110110111010011110110000000;
   assign mem[288159:288128] = 32'b00000000001011100001100110111011;
   assign mem[288191:288160] = 32'b00000111011110101000000100111000;
   assign mem[288223:288192] = 32'b00000011101001100110100010110100;
   assign mem[288255:288224] = 32'b11111001101010000001111111111000;
   assign mem[288287:288256] = 32'b00000010110111011101110011001000;
   assign mem[288319:288288] = 32'b11111100111100011111111011101100;
   assign mem[288351:288320] = 32'b00000110110000111001110001011000;
   assign mem[288383:288352] = 32'b11111000100011101110001100110000;
   assign mem[288415:288384] = 32'b00001000100001000100110100100000;
   assign mem[288447:288416] = 32'b11111000100100111111110111111000;
   assign mem[288479:288448] = 32'b00000010110101111001101010111000;
   assign mem[288511:288480] = 32'b11101100111101110110000110100000;
   assign mem[288543:288512] = 32'b11111111010001100010010011110010;
   assign mem[288575:288544] = 32'b00000011101101110010001100000000;
   assign mem[288607:288576] = 32'b00000101001100000110000000011000;
   assign mem[288639:288608] = 32'b00000000011001011000011110001111;
   assign mem[288671:288640] = 32'b11111101100111011101100011010100;
   assign mem[288703:288672] = 32'b00000000110111000011100010110010;
   assign mem[288735:288704] = 32'b00000000111101010010101001101011;
   assign mem[288767:288736] = 32'b00000111010000010001000111011000;
   assign mem[288799:288768] = 32'b00000010111100001000110001100100;
   assign mem[288831:288800] = 32'b11111010011011101010100100000000;
   assign mem[288863:288832] = 32'b11111011010011110110111000011000;
   assign mem[288895:288864] = 32'b00000001100000101100010011100000;
   assign mem[288927:288896] = 32'b00000100111000100110100011010000;
   assign mem[288959:288928] = 32'b00000000101010101111111101101001;
   assign mem[288991:288960] = 32'b00001000111101001110101101100000;
   assign mem[289023:288992] = 32'b11110110001110101111110001010000;
   assign mem[289055:289024] = 32'b00000110010001001110011101010000;
   assign mem[289087:289056] = 32'b11111111011101011011001100001000;
   assign mem[289119:289088] = 32'b00000111110001101000011001010000;
   assign mem[289151:289120] = 32'b11100101101010001101011110000000;
   assign mem[289183:289152] = 32'b11101100011101101100011101100000;
   assign mem[289215:289184] = 32'b00000011111110111011011011110000;
   assign mem[289247:289216] = 32'b00001001011011110010000111010000;
   assign mem[289279:289248] = 32'b00000000000000001101111101001100;
   assign mem[289311:289280] = 32'b11110010000000001000011100110000;
   assign mem[289343:289312] = 32'b00000001110001100100110100110000;
   assign mem[289375:289344] = 32'b00000001011100001101101111110100;
   assign mem[289407:289376] = 32'b00000110010011100100010101001000;
   assign mem[289439:289408] = 32'b11111000110010111001010111010000;
   assign mem[289471:289440] = 32'b00000100000100101000111100001000;
   assign mem[289503:289472] = 32'b00001000011100011011000000100000;
   assign mem[289535:289504] = 32'b00000001110000100000010111100100;
   assign mem[289567:289536] = 32'b11111100110111101001111001000100;
   assign mem[289599:289568] = 32'b11111000011001010000000111110000;
   assign mem[289631:289600] = 32'b00000000000101001100110011111000;
   assign mem[289663:289632] = 32'b11111111010101111010010000100011;
   assign mem[289695:289664] = 32'b00000000011010010000100111000110;
   assign mem[289727:289696] = 32'b00000000101000111000111001101110;
   assign mem[289759:289728] = 32'b11110010011111110100010000000000;
   assign mem[289791:289760] = 32'b11110111111010001110111110110000;
   assign mem[289823:289792] = 32'b11111001001011010101111001111000;
   assign mem[289855:289824] = 32'b00000100100111010001010100101000;
   assign mem[289887:289856] = 32'b00000100110111110111010100011000;
   assign mem[289919:289888] = 32'b11111110101010110000111010111110;
   assign mem[289951:289920] = 32'b00000001011011110101010101001010;
   assign mem[289983:289952] = 32'b11110001110011111000110011010000;
   assign mem[290015:289984] = 32'b00000100000110111010101100011000;
   assign mem[290047:290016] = 32'b11110100100101110000100100110000;
   assign mem[290079:290048] = 32'b00001011000010000100001101010000;
   assign mem[290111:290080] = 32'b11110100010100010011111100010000;
   assign mem[290143:290112] = 32'b00001001110110000111110111000000;
   assign mem[290175:290144] = 32'b00000010011110110111100010111000;
   assign mem[290207:290176] = 32'b00000011100111100110010011100000;
   assign mem[290239:290208] = 32'b11110000100000000011010001110000;
   assign mem[290271:290240] = 32'b00000101101010011110000101001000;
   assign mem[290303:290272] = 32'b00000010011010111000101101110000;
   assign mem[290335:290304] = 32'b11101111111111111111100111000000;
   assign mem[290367:290336] = 32'b00000011010011000101011010110000;
   assign mem[290399:290368] = 32'b00000001001100001110000110001100;
   assign mem[290431:290400] = 32'b00000101100101110011111101101000;
   assign mem[290463:290432] = 32'b00000100100001011101010110101000;
   assign mem[290495:290464] = 32'b11111101010101110101111000101100;
   assign mem[290527:290496] = 32'b00000010000100011100110110000100;
   assign mem[290559:290528] = 32'b11110011100111010111100101010000;
   assign mem[290591:290560] = 32'b11101111111100000010101011100000;
   assign mem[290623:290592] = 32'b11111011010000010011010001100000;
   assign mem[290655:290624] = 32'b00000100111011000001111000000000;
   assign mem[290687:290656] = 32'b00000010111001101010110100111000;
   assign mem[290719:290688] = 32'b00000101111100010010110101001000;
   assign mem[290751:290720] = 32'b00000000101100010111110111000000;
   assign mem[290783:290752] = 32'b11111111010011000111011111010110;
   assign mem[290815:290784] = 32'b00000101110110110110001011110000;
   assign mem[290847:290816] = 32'b11111111111111001101011000000100;
   assign mem[290879:290848] = 32'b11101010001101011100011011000000;
   assign mem[290911:290880] = 32'b11110110111000010011111011000000;
   assign mem[290943:290912] = 32'b11111100100111101110111101000100;
   assign mem[290975:290944] = 32'b00000000011101001100101110001110;
   assign mem[291007:290976] = 32'b00000110110000000011101011100000;
   assign mem[291039:291008] = 32'b00000010111101000001100111100100;
   assign mem[291071:291040] = 32'b00000100100001010100001101010000;
   assign mem[291103:291072] = 32'b00000010100001010001000011010100;
   assign mem[291135:291104] = 32'b00000011011001110010000101000100;
   assign mem[291167:291136] = 32'b00000010001111010111011101111100;
   assign mem[291199:291168] = 32'b11110101101000011001011100110000;
   assign mem[291231:291200] = 32'b11111010011110100111001100000000;
   assign mem[291263:291232] = 32'b11110110100011010010100111000000;
   assign mem[291295:291264] = 32'b00000010001111000111000000011000;
   assign mem[291327:291296] = 32'b00001000011101001110111010000000;
   assign mem[291359:291328] = 32'b00001001001010000000000110000000;
   assign mem[291391:291360] = 32'b11110111101110101011101001000000;
   assign mem[291423:291392] = 32'b11111010100010010110110001011000;
   assign mem[291455:291424] = 32'b00000011000100010101010100010100;
   assign mem[291487:291456] = 32'b00000010111100000100101100110100;
   assign mem[291519:291488] = 32'b11111011000010011011110001100000;
   assign mem[291551:291520] = 32'b00000111000101000001100011011000;
   assign mem[291583:291552] = 32'b11110011000001100110111101010000;
   assign mem[291615:291584] = 32'b00001000101000011001100100100000;
   assign mem[291647:291616] = 32'b11101011101111010001000101000000;
   assign mem[291679:291648] = 32'b11111010001100010101110001101000;
   assign mem[291711:291680] = 32'b11110011111000110101100001110000;
   assign mem[291743:291712] = 32'b11111111001111001001101000011000;
   assign mem[291775:291744] = 32'b00000010110100000010011001110000;
   assign mem[291807:291776] = 32'b00000100010011001000001010010000;
   assign mem[291839:291808] = 32'b11110010001110011011110101100000;
   assign mem[291871:291840] = 32'b11111100011010101101100011101100;
   assign mem[291903:291872] = 32'b00000000000010001110011101101110;
   assign mem[291935:291904] = 32'b00000111100100010011001001001000;
   assign mem[291967:291936] = 32'b11110001110110011010000010110000;
   assign mem[291999:291968] = 32'b00000100100100110001010100101000;
   assign mem[292031:292000] = 32'b00000000111111010100011101110110;
   assign mem[292063:292032] = 32'b11111001111011111100111010111000;
   assign mem[292095:292064] = 32'b00000000100000010100110111111101;
   assign mem[292127:292096] = 32'b00001000110001100011001111000000;
   assign mem[292159:292128] = 32'b11111101011111110000011011001000;
   assign mem[292191:292160] = 32'b00000111000011000100000110010000;
   assign mem[292223:292192] = 32'b11111100101011100001101000011000;
   assign mem[292255:292224] = 32'b11111001001001111001011000101000;
   assign mem[292287:292256] = 32'b00000010001101110111110011111000;
   assign mem[292319:292288] = 32'b11111101011100001100100101100000;
   assign mem[292351:292320] = 32'b11111111101010000011001001101000;
   assign mem[292383:292352] = 32'b00000101010011101100011001011000;
   assign mem[292415:292384] = 32'b11111111100101011000001001010100;
   assign mem[292447:292416] = 32'b00000001000001001011110111010100;
   assign mem[292479:292448] = 32'b11111111001101111011000000111101;
   assign mem[292511:292480] = 32'b11101011011111011101111010000000;
   assign mem[292543:292512] = 32'b11110011001100010100101000010000;
   assign mem[292575:292544] = 32'b11110110001000001101001110000000;
   assign mem[292607:292576] = 32'b00000110110001111001010010000000;
   assign mem[292639:292608] = 32'b00000000000000010000110110011001;
   assign mem[292671:292640] = 32'b00000111011110011001010000101000;
   assign mem[292703:292672] = 32'b00000100001110001111010100000000;
   assign mem[292735:292704] = 32'b11111110001000101011010000011100;
   assign mem[292767:292736] = 32'b00000011110000001001000011111000;
   assign mem[292799:292768] = 32'b11111110001000011011110110000000;
   assign mem[292831:292800] = 32'b00000010110110100011001110010100;
   assign mem[292863:292832] = 32'b11100011010000110111010110000000;
   assign mem[292895:292864] = 32'b11111111110000100000001100001110;
   assign mem[292927:292896] = 32'b00000101001111000111011111011000;
   assign mem[292959:292928] = 32'b00000000010010001001000101111000;
   assign mem[292991:292960] = 32'b11111111001101111011010011111101;
   assign mem[293023:292992] = 32'b00000100111001100011011000011000;
   assign mem[293055:293024] = 32'b11111100000000000001011111010000;
   assign mem[293087:293056] = 32'b00000110011100001101011101101000;
   assign mem[293119:293088] = 32'b11111010010001110101010001010000;
   assign mem[293151:293120] = 32'b00001001001010000110011011000000;
   assign mem[293183:293152] = 32'b11111100101100110111001010100100;
   assign mem[293215:293184] = 32'b11111111010011100000110110110101;
   assign mem[293247:293216] = 32'b11101011001111101011010110000000;
   assign mem[293279:293248] = 32'b00001101001111101010011001000000;
   assign mem[293311:293280] = 32'b11110000011111000100000100000000;
   assign mem[293343:293312] = 32'b11111100000110011010000111111000;
   assign mem[293375:293344] = 32'b00001110101101101011010111010000;
   assign mem[293407:293376] = 32'b11101111010110010011001101100000;
   assign mem[293439:293408] = 32'b11111010001010001100111100110000;
   assign mem[293471:293440] = 32'b11111011001010110101001101000000;
   assign mem[293503:293472] = 32'b11110110000001111101010010110000;
   assign mem[293535:293504] = 32'b00000111101010001010001111000000;
   assign mem[293567:293536] = 32'b11111100001101010000011001111100;
   assign mem[293599:293568] = 32'b00000001100111111001011111101110;
   assign mem[293631:293600] = 32'b11111111110000101010111111100001;
   assign mem[293663:293632] = 32'b00000101000001110111100010101000;
   assign mem[293695:293664] = 32'b11111001110000101100110010010000;
   assign mem[293727:293696] = 32'b00000101010010000110001110000000;
   assign mem[293759:293728] = 32'b11111001101101110001001010111000;
   assign mem[293791:293760] = 32'b00000011110100010100111000101100;
   assign mem[293823:293792] = 32'b11111000110010001010100010011000;
   assign mem[293855:293824] = 32'b00000111010010111001101010011000;
   assign mem[293887:293856] = 32'b00000001100101101111101110011000;
   assign mem[293919:293888] = 32'b00000000101011000100011110101110;
   assign mem[293951:293920] = 32'b11101111011101010101101101100000;
   assign mem[293983:293952] = 32'b11110101111101001010001111010000;
   assign mem[294015:293984] = 32'b00000011101000001000100011111100;
   assign mem[294047:294016] = 32'b00001000111000101101100000110000;
   assign mem[294079:294048] = 32'b11111110100100010011011000000110;
   assign mem[294111:294080] = 32'b00000010001110111011110111111000;
   assign mem[294143:294112] = 32'b11111100110010110011101001011000;
   assign mem[294175:294144] = 32'b11111010001101110001100001110000;
   assign mem[294207:294176] = 32'b00000011001001110011101110001000;
   assign mem[294239:294208] = 32'b00000111111111101010101001001000;
   assign mem[294271:294240] = 32'b00000010111010011010001000001000;
   assign mem[294303:294272] = 32'b11111110011101000000001111010100;
   assign mem[294335:294304] = 32'b11111110101101110110010110000000;
   assign mem[294367:294336] = 32'b11111110111010000100010100101100;
   assign mem[294399:294368] = 32'b00000100100110001100010101110000;
   assign mem[294431:294400] = 32'b00000100100101110100011000100000;
   assign mem[294463:294432] = 32'b00000000111101101100001101011011;
   assign mem[294495:294464] = 32'b11111111001100100100110101010000;
   assign mem[294527:294496] = 32'b11111111101110010000111001000011;
   assign mem[294559:294528] = 32'b00000101000110111111011011001000;
   assign mem[294591:294560] = 32'b11111111001010110000011010011010;
   assign mem[294623:294592] = 32'b11111010011111010110110110110000;
   assign mem[294655:294624] = 32'b00000010000111101100101111101100;
   assign mem[294687:294656] = 32'b11111000011100011010000110010000;
   assign mem[294719:294688] = 32'b11111111100101011001101011010101;
   assign mem[294751:294720] = 32'b11111100101011010100101101011100;
   assign mem[294783:294752] = 32'b00000001010000111010000100011010;
   assign mem[294815:294784] = 32'b00000000001010111111100011101011;
   assign mem[294847:294816] = 32'b00000010011011101111001111011100;
   assign mem[294879:294848] = 32'b00000010010110011101101110010000;
   assign mem[294911:294880] = 32'b11111110011111010101000011100100;
   assign mem[294943:294912] = 32'b11111010101100101110010001111000;
   assign mem[294975:294944] = 32'b00000000000101011001011111001001;
   assign mem[295007:294976] = 32'b11111101000001110110110001100100;
   assign mem[295039:295008] = 32'b00000010110111001100010100011000;
   assign mem[295071:295040] = 32'b11111111000100101100000101001101;
   assign mem[295103:295072] = 32'b00000010000000011001010110111000;
   assign mem[295135:295104] = 32'b00000000101110010110011111011100;
   assign mem[295167:295136] = 32'b00000001100110001101101000110010;
   assign mem[295199:295168] = 32'b00000000110000001101111110100000;
   assign mem[295231:295200] = 32'b11111100001011111001101010101000;
   assign mem[295263:295232] = 32'b11110101101000010011100110110000;
   assign mem[295295:295264] = 32'b00000010000011111110001011100100;
   assign mem[295327:295296] = 32'b11111110101000100101100101100000;
   assign mem[295359:295328] = 32'b11111110111011100101001110110100;
   assign mem[295391:295360] = 32'b11110111011101000001101100100000;
   assign mem[295423:295392] = 32'b00000100101010011011000001100000;
   assign mem[295455:295424] = 32'b00000111110100010011100000010000;
   assign mem[295487:295456] = 32'b00000001100111101010111110001110;
   assign mem[295519:295488] = 32'b11111010111100111010010001110000;
   assign mem[295551:295520] = 32'b11110111101011001011110101100000;
   assign mem[295583:295552] = 32'b11110010000111010100101001100000;
   assign mem[295615:295584] = 32'b11111111011100111010000001000111;
   assign mem[295647:295616] = 32'b00001000010100111100001001110000;
   assign mem[295679:295648] = 32'b00000110111001000110110010001000;
   assign mem[295711:295680] = 32'b11111101000100100001011110110000;
   assign mem[295743:295712] = 32'b11111000101100000111101100101000;
   assign mem[295775:295744] = 32'b00000010000010111001110000010100;
   assign mem[295807:295776] = 32'b00001000001110110110100110110000;
   assign mem[295839:295808] = 32'b00000010001111111001111000011100;
   assign mem[295871:295840] = 32'b11101101011001000111011100100000;
   assign mem[295903:295872] = 32'b00000000100110001001010110001000;
   assign mem[295935:295904] = 32'b00001000001111101001110100100000;
   assign mem[295967:295936] = 32'b00000100000110110010101111001000;
   assign mem[295999:295968] = 32'b11110101010011111111000010010000;
   assign mem[296031:296000] = 32'b11110111000010000111110100000000;
   assign mem[296063:296032] = 32'b00000001100001000001010100000000;
   assign mem[296095:296064] = 32'b00000011010101010000001011100000;
   assign mem[296127:296096] = 32'b00000101100100111011100110010000;
   assign mem[296159:296128] = 32'b11110101101111110000100011000000;
   assign mem[296191:296160] = 32'b00000011001011110001010101010100;
   assign mem[296223:296192] = 32'b00001010000010101110011001000000;
   assign mem[296255:296224] = 32'b11111110110110001011001100011100;
   assign mem[296287:296256] = 32'b11111011001100101000110100000000;
   assign mem[296319:296288] = 32'b11110100000100001111110001110000;
   assign mem[296351:296320] = 32'b00000010100011100111001000101000;
   assign mem[296383:296352] = 32'b11111011111100001011001101010000;
   assign mem[296415:296384] = 32'b00000010111110111111111000001100;
   assign mem[296447:296416] = 32'b11110111011100111001010100010000;
   assign mem[296479:296448] = 32'b00000101011000011010000111010000;
   assign mem[296511:296480] = 32'b11111101111011110111110101100100;
   assign mem[296543:296512] = 32'b11111000110101110101110111101000;
   assign mem[296575:296544] = 32'b00000000001111011001001111001100;
   assign mem[296607:296576] = 32'b11111100111111110101100010110100;
   assign mem[296639:296608] = 32'b00000010000010001101101110001000;
   assign mem[296671:296640] = 32'b00000001101100110101111100010000;
   assign mem[296703:296672] = 32'b11111101110111110110001011100000;
   assign mem[296735:296704] = 32'b11111111010100111011110001010001;
   assign mem[296767:296736] = 32'b11110101110100011111001111000000;
   assign mem[296799:296768] = 32'b00000101001100010001001101110000;
   assign mem[296831:296800] = 32'b00000010100100011111100010111000;
   assign mem[296863:296832] = 32'b11111000001011101010110001111000;
   assign mem[296895:296864] = 32'b11111111111010011110111110000100;
   assign mem[296927:296896] = 32'b00000001101011001010110001011010;
   assign mem[296959:296928] = 32'b11111110111010010000000011000000;
   assign mem[296991:296960] = 32'b11111110100111110100100011110100;
   assign mem[297023:296992] = 32'b11110111111011110101011100000000;
   assign mem[297055:297024] = 32'b11111111111111001011001010001101;
   assign mem[297087:297056] = 32'b00000001010000000001111111111000;
   assign mem[297119:297088] = 32'b11111110100110011110101111110010;
   assign mem[297151:297120] = 32'b11101100010100111111001100100000;
   assign mem[297183:297152] = 32'b11111100010111001111001010100000;
   assign mem[297215:297184] = 32'b00000000000100010110000110100101;
   assign mem[297247:297216] = 32'b00001011101101000111110011010000;
   assign mem[297279:297248] = 32'b11111110110011111101101010001100;
   assign mem[297311:297280] = 32'b00001001111100101010000100100000;
   assign mem[297343:297312] = 32'b11111010100110110111111010001000;
   assign mem[297375:297344] = 32'b11111100100110010000110100100100;
   assign mem[297407:297376] = 32'b11110000010100111111001011100000;
   assign mem[297439:297408] = 32'b00001000000101010000111001110000;
   assign mem[297471:297440] = 32'b11110101110111101011101011110000;
   assign mem[297503:297472] = 32'b11111110010011010110111010011100;
   assign mem[297535:297504] = 32'b00000011011100000101001110110100;
   assign mem[297567:297536] = 32'b11111110001011010101001001010110;
   assign mem[297599:297568] = 32'b11111000011010101111100110011000;
   assign mem[297631:297600] = 32'b11111110010010000101001101001000;
   assign mem[297663:297632] = 32'b00000011001100110110110010101100;
   assign mem[297695:297664] = 32'b00000111001000110100110011110000;
   assign mem[297727:297696] = 32'b11110100101100000101011001100000;
   assign mem[297759:297728] = 32'b00000111010100101010001000001000;
   assign mem[297791:297760] = 32'b11111000100010100011001010011000;
   assign mem[297823:297792] = 32'b00000010011001100001101100110100;
   assign mem[297855:297824] = 32'b00000100001011111000000000100000;
   assign mem[297887:297856] = 32'b00000001010111110100010010111010;
   assign mem[297919:297888] = 32'b11111010010101000100100100100000;
   assign mem[297951:297920] = 32'b00000010001011011111001000101100;
   assign mem[297983:297952] = 32'b11111110011010011100100111000110;
   assign mem[298015:297984] = 32'b00000000000111000001110010001001;
   assign mem[298047:298016] = 32'b00000010110010001011100100110100;
   assign mem[298079:298048] = 32'b00000000010110100010011011000010;
   assign mem[298111:298080] = 32'b11101110000011011000100110000000;
   assign mem[298143:298112] = 32'b11110101100010001100010001000000;
   assign mem[298175:298144] = 32'b00000011100010100011010000010100;
   assign mem[298207:298176] = 32'b00000011110000100101011101101000;
   assign mem[298239:298208] = 32'b00000010000001010100011000000100;
   assign mem[298271:298240] = 32'b11111000100111011111110010110000;
   assign mem[298303:298272] = 32'b11110100101000010100010101100000;
   assign mem[298335:298304] = 32'b11111010011011100110010011010000;
   assign mem[298367:298336] = 32'b00000101001101010111000100001000;
   assign mem[298399:298368] = 32'b11111000111000101010011100011000;
   assign mem[298431:298400] = 32'b00000011010100000110001100000100;
   assign mem[298463:298432] = 32'b00000101111010101100010001000000;
   assign mem[298495:298464] = 32'b11111011100110001110100000000000;
   assign mem[298527:298496] = 32'b00000010000110110101000111111100;
   assign mem[298559:298528] = 32'b00000001001100100110001011111100;
   assign mem[298591:298560] = 32'b00000001111100010001010011010010;
   assign mem[298623:298592] = 32'b11110011010100010101110100010000;
   assign mem[298655:298624] = 32'b11111000001010011001111001111000;
   assign mem[298687:298656] = 32'b00000010100110110010001000011000;
   assign mem[298719:298688] = 32'b00000001000001101001010111011000;
   assign mem[298751:298720] = 32'b00000000101101011110111110100111;
   assign mem[298783:298752] = 32'b00000111100000101100110010111000;
   assign mem[298815:298784] = 32'b11111111000111000101101111101000;
   assign mem[298847:298816] = 32'b11111101110110110010100110110000;
   assign mem[298879:298848] = 32'b00000010110100101000110011010100;
   assign mem[298911:298880] = 32'b11111100100100100100000110000000;
   assign mem[298943:298912] = 32'b11111101011110000101001110000000;
   assign mem[298975:298944] = 32'b00000111100011111110000001101000;
   assign mem[299007:298976] = 32'b11110111011100100101110111110000;
   assign mem[299039:299008] = 32'b00001100110110110100110010110000;
   assign mem[299071:299040] = 32'b11111011111110010010111010011000;
   assign mem[299103:299072] = 32'b11110110100010100110101010100000;
   assign mem[299135:299104] = 32'b00000110110101010110110011010000;
   assign mem[299167:299136] = 32'b11111111100001010011111010110000;
   assign mem[299199:299168] = 32'b11111101000011101111010001100000;
   assign mem[299231:299200] = 32'b00000110101110000101100001000000;
   assign mem[299263:299232] = 32'b00000011011010001001000100001000;
   assign mem[299295:299264] = 32'b00000110001010111000111111011000;
   assign mem[299327:299296] = 32'b11111000111011101100011101110000;
   assign mem[299359:299328] = 32'b11101011010000101101010000000000;
   assign mem[299391:299360] = 32'b00001000101000110011011000110000;
   assign mem[299423:299392] = 32'b00000011000110101101000010110000;
   assign mem[299455:299424] = 32'b11101110001111000010111011000000;
   assign mem[299487:299456] = 32'b11111001101100001010110011110000;
   assign mem[299519:299488] = 32'b11110110100010000100100001110000;
   assign mem[299551:299520] = 32'b00000110010101101100100000110000;
   assign mem[299583:299552] = 32'b00000001101100110101111000100010;
   assign mem[299615:299584] = 32'b11111010111010010100010010010000;
   assign mem[299647:299616] = 32'b11111011111111000111101011011000;
   assign mem[299679:299648] = 32'b00000100110100110101000001100000;
   assign mem[299711:299680] = 32'b00000101100001101010010101101000;
   assign mem[299743:299712] = 32'b11111101100100111101011010001000;
   assign mem[299775:299744] = 32'b00001000110000101010011001010000;
   assign mem[299807:299776] = 32'b00000000000011011011100111111011;
   assign mem[299839:299808] = 32'b11111010101100111111000101110000;
   assign mem[299871:299840] = 32'b11110001011011110000101001100000;
   assign mem[299903:299872] = 32'b11111101101011110101100010000100;
   assign mem[299935:299904] = 32'b11110111011110101111101101000000;
   assign mem[299967:299936] = 32'b00000101000001001101000011111000;
   assign mem[299999:299968] = 32'b00000010111011111111000011001000;
   assign mem[300031:300000] = 32'b11111111011111101010100011000100;
   assign mem[300063:300032] = 32'b11111011101010010001111110010000;
   assign mem[300095:300064] = 32'b11111011101111110010111100100000;
   assign mem[300127:300096] = 32'b11111110011101001111011110100000;
   assign mem[300159:300128] = 32'b00000110001001111111110110111000;
   assign mem[300191:300160] = 32'b00000011111001000110011001000100;
   assign mem[300223:300192] = 32'b00001011111100001110000000010000;
   assign mem[300255:300224] = 32'b11110111010100110111010011100000;
   assign mem[300287:300256] = 32'b11111001000111010110110010010000;
   assign mem[300319:300288] = 32'b11111001100110111011101001000000;
   assign mem[300351:300320] = 32'b00001111111010110101100011000000;
   assign mem[300383:300352] = 32'b00000000101000101111011101110011;
   assign mem[300415:300384] = 32'b11110000110110000100010001100000;
   assign mem[300447:300416] = 32'b11111010010000101111001111011000;
   assign mem[300479:300448] = 32'b11111111110110011100101111000001;
   assign mem[300511:300480] = 32'b00000001001010000001100111011110;
   assign mem[300543:300512] = 32'b11111101100011110011001010101000;
   assign mem[300575:300544] = 32'b11111111001100101100011000010010;
   assign mem[300607:300576] = 32'b00000010000101101101001101000100;
   assign mem[300639:300608] = 32'b00000010110001101001100111011000;
   assign mem[300671:300640] = 32'b11111111100011001111101110110011;
   assign mem[300703:300672] = 32'b00000011011011101100001110010000;
   assign mem[300735:300704] = 32'b11111101101111110101010011000000;
   assign mem[300767:300736] = 32'b11111101001100110111110100111000;
   assign mem[300799:300768] = 32'b00000010100111111111101111111000;
   assign mem[300831:300800] = 32'b00001011001000011101001001000000;
   assign mem[300863:300832] = 32'b11111010010111000000110001000000;
   assign mem[300895:300864] = 32'b11111111101110011110000000111001;
   assign mem[300927:300896] = 32'b00000011100111110110000110110100;
   assign mem[300959:300928] = 32'b00000101100010100110110001111000;
   assign mem[300991:300960] = 32'b11111001110101101110110111011000;
   assign mem[301023:300992] = 32'b11111011010101110101111011111000;
   assign mem[301055:301024] = 32'b00000011110101001100010011100000;
   assign mem[301087:301056] = 32'b11111010111001001101001010101000;
   assign mem[301119:301088] = 32'b00000011111010000000111010101100;
   assign mem[301151:301120] = 32'b00000011111111110011100111110000;
   assign mem[301183:301152] = 32'b11110001000001100110110000000000;
   assign mem[301215:301184] = 32'b11111011101010110000010001010000;
   assign mem[301247:301216] = 32'b00000000010001111100111100110100;
   assign mem[301279:301248] = 32'b11110101101110001011011001000000;
   assign mem[301311:301280] = 32'b00000100100101101000111000011000;
   assign mem[301343:301312] = 32'b00000101001101010011000100101000;
   assign mem[301375:301344] = 32'b00000000001011110111011110110011;
   assign mem[301407:301376] = 32'b00000000110100001110011101011000;
   assign mem[301439:301408] = 32'b00000001110001001101011010100010;
   assign mem[301471:301440] = 32'b00001010101101001100100011000000;
   assign mem[301503:301472] = 32'b11111110100010111111011100101110;
   assign mem[301535:301504] = 32'b11110010110110101000111011100000;
   assign mem[301567:301536] = 32'b11111000010111100001111100110000;
   assign mem[301599:301568] = 32'b11110101100111010101110101110000;
   assign mem[301631:301600] = 32'b00001001010110100000101001110000;
   assign mem[301663:301632] = 32'b00000000111011011111101001101100;
   assign mem[301695:301664] = 32'b00001011111011100010011111000000;
   assign mem[301727:301696] = 32'b11111001100000000100101110100000;
   assign mem[301759:301728] = 32'b11100100101100111100010011100000;
   assign mem[301791:301760] = 32'b11111111101110101000110111011000;
   assign mem[301823:301792] = 32'b11111110010110010010101001011000;
   assign mem[301855:301824] = 32'b11111110100011010010000001100000;
   assign mem[301887:301856] = 32'b00000010100101101011001011110100;
   assign mem[301919:301888] = 32'b00000001100000110101000000111000;
   assign mem[301951:301920] = 32'b11111101111111010111000000011100;
   assign mem[301983:301952] = 32'b11111011011111000000010011110000;
   assign mem[302015:301984] = 32'b00000000110111010010110101100010;
   assign mem[302047:302016] = 32'b11111101000000110010111110001100;
   assign mem[302079:302048] = 32'b11111011111110001010110100111000;
   assign mem[302111:302080] = 32'b11111100010010011000100101001000;
   assign mem[302143:302112] = 32'b11111101100101000101100100111000;
   assign mem[302175:302144] = 32'b11111001010001111101100011100000;
   assign mem[302207:302176] = 32'b11111011111100010010100010100000;
   assign mem[302239:302208] = 32'b00000011101011000010011000110000;
   assign mem[302271:302240] = 32'b11110111110010001010100110010000;
   assign mem[302303:302272] = 32'b00000011010011100011101100001100;
   assign mem[302335:302304] = 32'b00001000000011101110000010000000;
   assign mem[302367:302336] = 32'b11111011111100101111110011101000;
   assign mem[302399:302368] = 32'b00000101001110001010111101110000;
   assign mem[302431:302400] = 32'b00000000101100001100010110111010;
   assign mem[302463:302432] = 32'b11111101101000000101001111110000;
   assign mem[302495:302464] = 32'b00001101111101011110111110100000;
   assign mem[302527:302496] = 32'b11110010110101000001110000100000;
   assign mem[302559:302528] = 32'b00000001010100101000111110001010;
   assign mem[302591:302560] = 32'b11110100010010001101010010100000;
   assign mem[302623:302592] = 32'b11111010100111011110101110100000;
   assign mem[302655:302624] = 32'b11110100011101110100111111000000;
   assign mem[302687:302656] = 32'b00001000100110011010010111000000;
   assign mem[302719:302688] = 32'b11111001001010001001000011001000;
   assign mem[302751:302720] = 32'b00000010001000000101011100000000;
   assign mem[302783:302752] = 32'b11110011011000000100000100000000;
   assign mem[302815:302784] = 32'b00000110111011111100110110100000;
   assign mem[302847:302816] = 32'b11111001000111100011110110001000;
   assign mem[302879:302848] = 32'b11111101111010111111001011101100;
   assign mem[302911:302880] = 32'b11101100010011010000100111100000;
   assign mem[302943:302912] = 32'b00000010101100001110011001011100;
   assign mem[302975:302944] = 32'b00000010111010101000101001001100;
   assign mem[303007:302976] = 32'b00001011100111100101101011000000;
   assign mem[303039:303008] = 32'b00000001001011010111111110000100;
   assign mem[303071:303040] = 32'b00010000001011101111111011000000;
   assign mem[303103:303072] = 32'b00000111100011011000010111101000;
   assign mem[303135:303104] = 32'b11111111001010001100011111011100;
   assign mem[303167:303136] = 32'b11101011011010000011101011100000;
   assign mem[303199:303168] = 32'b11110010111100101111010110100000;
   assign mem[303231:303200] = 32'b11111011011011100001111011101000;
   assign mem[303263:303232] = 32'b11111100110001001011011110111100;
   assign mem[303295:303264] = 32'b00000000001100011000000000000011;
   assign mem[303327:303296] = 32'b11111100100110000001000000011000;
   assign mem[303359:303328] = 32'b11111100000011000101001010101100;
   assign mem[303391:303360] = 32'b00000010001011101111000100111000;
   assign mem[303423:303392] = 32'b11110100100011010100000101000000;
   assign mem[303455:303424] = 32'b00000101100010101001111101000000;
   assign mem[303487:303456] = 32'b11111010010111011010000011110000;
   assign mem[303519:303488] = 32'b00000000100101010110101000100100;
   assign mem[303551:303520] = 32'b00000000111000111110111001110110;
   assign mem[303583:303552] = 32'b11111100011111111100000101011100;
   assign mem[303615:303584] = 32'b00000011111100101010101110010100;
   assign mem[303647:303616] = 32'b00000111111100111110110100111000;
   assign mem[303679:303648] = 32'b11110110000111001110001111100000;
   assign mem[303711:303680] = 32'b11110110011100111111110101110000;
   assign mem[303743:303712] = 32'b11110000010011111000011001010000;
   assign mem[303775:303744] = 32'b00000010111010011011101001111100;
   assign mem[303807:303776] = 32'b00000001000100000100111001010100;
   assign mem[303839:303808] = 32'b00000010011000100010011111110000;
   assign mem[303871:303840] = 32'b00000111011111111011100100101000;
   assign mem[303903:303872] = 32'b00000001010100111100000100111100;
   assign mem[303935:303904] = 32'b00000001011101010001001111000000;
   assign mem[303967:303936] = 32'b00000000010101000001101110101101;
   assign mem[303999:303968] = 32'b11110001100110100111111010010000;
   assign mem[304031:304000] = 32'b11111110101100111101101011011100;
   assign mem[304063:304032] = 32'b11111101011011100100110111110000;
   assign mem[304095:304064] = 32'b00000100011010000010001000101000;
   assign mem[304127:304096] = 32'b11111011011000101010011000011000;
   assign mem[304159:304128] = 32'b00000111011011001100000110010000;
   assign mem[304191:304160] = 32'b11111001010110110000110111111000;
   assign mem[304223:304192] = 32'b11110101010010011011100010110000;
   assign mem[304255:304224] = 32'b11111100011110100100100010000000;
   assign mem[304287:304256] = 32'b00001101000111100110010000010000;
   assign mem[304319:304288] = 32'b00000101110000111010000011101000;
   assign mem[304351:304320] = 32'b11111111111000010011001101111111;
   assign mem[304383:304352] = 32'b11110111100101011000111100110000;
   assign mem[304415:304384] = 32'b00000010101011101111010100000000;
   assign mem[304447:304416] = 32'b00000011011110001111100000100100;
   assign mem[304479:304448] = 32'b00000000101110001011010111001010;
   assign mem[304511:304480] = 32'b11111011010100101011101011101000;
   assign mem[304543:304512] = 32'b11110101101000110011110111010000;
   assign mem[304575:304544] = 32'b00000100000001011101001101000000;
   assign mem[304607:304576] = 32'b00000010000111110011101110100000;
   assign mem[304639:304608] = 32'b00000010011000000111110011100000;
   assign mem[304671:304640] = 32'b11111101011111011001001000110000;
   assign mem[304703:304672] = 32'b11111000011100111001011100111000;
   assign mem[304735:304704] = 32'b11111100100111011101100001100000;
   assign mem[304767:304736] = 32'b00000110011010111111001101111000;
   assign mem[304799:304768] = 32'b00000000101110110100011100001101;
   assign mem[304831:304800] = 32'b11111110111110001100101101110010;
   assign mem[304863:304832] = 32'b00000110010001010011011011011000;
   assign mem[304895:304864] = 32'b00000010011001111101101100100000;
   assign mem[304927:304896] = 32'b11111000111011100001010111010000;
   assign mem[304959:304928] = 32'b00000111000001011100111100100000;
   assign mem[304991:304960] = 32'b00000110011111001110010010111000;
   assign mem[305023:304992] = 32'b00000011100001100111101001110000;
   assign mem[305055:305024] = 32'b11110110001000101100001100010000;
   assign mem[305087:305056] = 32'b11111001010011010010010111000000;
   assign mem[305119:305088] = 32'b11110101011011000100101000000000;
   assign mem[305151:305120] = 32'b00001000010111100101111110000000;
   assign mem[305183:305152] = 32'b00000011001010011000111101001000;
   assign mem[305215:305184] = 32'b11111110110000011110011011100010;
   assign mem[305247:305216] = 32'b00000001101011111001110110000110;
   assign mem[305279:305248] = 32'b11111010101110001001010010010000;
   assign mem[305311:305280] = 32'b11111001000001101111100011110000;
   assign mem[305343:305312] = 32'b00000000110010001000110111011110;
   assign mem[305375:305344] = 32'b11111110100110001001011110000110;
   assign mem[305407:305376] = 32'b11111111010110011100101100101110;
   assign mem[305439:305408] = 32'b11111110001110000001010110001110;
   assign mem[305471:305440] = 32'b00000011000100011111000110110100;
   assign mem[305503:305472] = 32'b00000100001100011110000101111000;
   assign mem[305535:305504] = 32'b00000010000110010101001000111000;
   assign mem[305567:305536] = 32'b11110111111111011110101010010000;
   assign mem[305599:305568] = 32'b00000010100111011010111011001100;
   assign mem[305631:305600] = 32'b11111111100010000000101011111011;
   assign mem[305663:305632] = 32'b11111110010101000010011110000110;
   assign mem[305695:305664] = 32'b11111110100010000001001101011010;
   assign mem[305727:305696] = 32'b00000000000010110110001100110101;
   assign mem[305759:305728] = 32'b00000001101010100110001001100000;
   assign mem[305791:305760] = 32'b00000101110000011110110101111000;
   assign mem[305823:305792] = 32'b00000101001111111001011101111000;
   assign mem[305855:305824] = 32'b11111011010100110110110010000000;
   assign mem[305887:305856] = 32'b11110111111010100101101010000000;
   assign mem[305919:305888] = 32'b11111111010010110110001001101110;
   assign mem[305951:305920] = 32'b11111101110010011011110111100100;
   assign mem[305983:305952] = 32'b00000011001001001011110001101100;
   assign mem[306015:305984] = 32'b00001100000001101000110001010000;
   assign mem[306047:306016] = 32'b11110101000010010111110001110000;
   assign mem[306079:306048] = 32'b11111100011010001101011010010000;
   assign mem[306111:306080] = 32'b11111010001000010111111111101000;
   assign mem[306143:306112] = 32'b00000000011111111110001110101010;
   assign mem[306175:306144] = 32'b11110110111111101001111100010000;
   assign mem[306207:306176] = 32'b11111001110011101010000111000000;
   assign mem[306239:306208] = 32'b00000101111111010101100110110000;
   assign mem[306271:306240] = 32'b00000000000110011111100011000100;
   assign mem[306303:306272] = 32'b11111011010001101001000110110000;
   assign mem[306335:306304] = 32'b00000010111000100111110100000100;
   assign mem[306367:306336] = 32'b11110001010000001011110110010000;
   assign mem[306399:306368] = 32'b11111111111111100110010000001110;
   assign mem[306431:306400] = 32'b11110100001110001000101110010000;
   assign mem[306463:306432] = 32'b11111001011101110110110110100000;
   assign mem[306495:306464] = 32'b00000000001101101101100101000100;
   assign mem[306527:306496] = 32'b00000000111010011001110001011110;
   assign mem[306559:306528] = 32'b00000000100011010101111001101000;
   assign mem[306591:306560] = 32'b00001011011110011111011010100000;
   assign mem[306623:306592] = 32'b11111001011111010110100100010000;
   assign mem[306655:306624] = 32'b00001101101111001001101001100000;
   assign mem[306687:306656] = 32'b11100110011000111010110100000000;
   assign mem[306719:306688] = 32'b00001100001011101100011001010000;
   assign mem[306751:306720] = 32'b11110001100100101101111111010000;
   assign mem[306783:306752] = 32'b11110010001100100000101101010000;
   assign mem[306815:306784] = 32'b11111001011101000010000011000000;
   assign mem[306847:306816] = 32'b11110010011011010001110000110000;
   assign mem[306879:306848] = 32'b11111011010001000110101000010000;
   assign mem[306911:306880] = 32'b00000100000110010111110101101000;
   assign mem[306943:306912] = 32'b11110111101100000001101101110000;
   assign mem[306975:306944] = 32'b00001000101010111111111000000000;
   assign mem[307007:306976] = 32'b11101001000011011001111111000000;
   assign mem[307039:307008] = 32'b00000100110000101111000100101000;
   assign mem[307071:307040] = 32'b11110100011010001111001000100000;
   assign mem[307103:307072] = 32'b11111011111011000101011001100000;
   assign mem[307135:307104] = 32'b00000010011101001000000010110100;
   assign mem[307167:307136] = 32'b11111110000001100111101101011010;
   assign mem[307199:307168] = 32'b11111101000000111011111100101100;
   assign mem[307231:307200] = 32'b11111010101101110111000011000000;
   assign mem[307263:307232] = 32'b00001010001000110101000100000000;
   assign mem[307295:307264] = 32'b00000100001001011110101000100000;
   assign mem[307327:307296] = 32'b00000011011001101101110110000100;
   assign mem[307359:307328] = 32'b00000010000010101101101111111000;
   assign mem[307391:307360] = 32'b11111111101101001111001011111000;
   assign mem[307423:307392] = 32'b11111010111110001100100010110000;
   assign mem[307455:307424] = 32'b11111010000110011110110001101000;
   assign mem[307487:307456] = 32'b11111010000000111110011100010000;
   assign mem[307519:307488] = 32'b00000110000110001000011011111000;
   assign mem[307551:307520] = 32'b11111010101001101011111000100000;
   assign mem[307583:307552] = 32'b11111101101011010100101010100100;
   assign mem[307615:307584] = 32'b11111001000101000101010111111000;
   assign mem[307647:307616] = 32'b00001010100100100011011101000000;
   assign mem[307679:307648] = 32'b11111110000110011110101101011010;
   assign mem[307711:307680] = 32'b11111111001111011110101101010010;
   assign mem[307743:307712] = 32'b00000100110001011101111111110000;
   assign mem[307775:307744] = 32'b00000011101010111101010100111000;
   assign mem[307807:307776] = 32'b11111100100100011011110010000000;
   assign mem[307839:307808] = 32'b11111011101001111011001100000000;
   assign mem[307871:307840] = 32'b11111100001111010111100111100000;
   assign mem[307903:307872] = 32'b11101101010110010111011001000000;
   assign mem[307935:307904] = 32'b11110100111110011101000100000000;
   assign mem[307967:307936] = 32'b00000011011000111100011111111000;
   assign mem[307999:307968] = 32'b00000101001000001101001110010000;
   assign mem[308031:308000] = 32'b00000010111110011011111110110000;
   assign mem[308063:308032] = 32'b00000001111011001001001000101100;
   assign mem[308095:308064] = 32'b11110000101111000011110000110000;
   assign mem[308127:308096] = 32'b11111011100100011011111011111000;
   assign mem[308159:308128] = 32'b11111100111111101011010010110100;
   assign mem[308191:308160] = 32'b11111111000011001101010100110001;
   assign mem[308223:308192] = 32'b00000110110000100100101110101000;
   assign mem[308255:308224] = 32'b11110101000011100011111010110000;
   assign mem[308287:308256] = 32'b00000000110110000100101111011001;
   assign mem[308319:308288] = 32'b00001000011101011101111110110000;
   assign mem[308351:308320] = 32'b00000010111011111010100001110100;
   assign mem[308383:308352] = 32'b11110111000001011111101010000000;
   assign mem[308415:308384] = 32'b11111011010100101010101111101000;
   assign mem[308447:308416] = 32'b11110111110000000111110101100000;
   assign mem[308479:308448] = 32'b00000000011010111100001010111011;
   assign mem[308511:308480] = 32'b11110001100101011010001001110000;
   assign mem[308543:308512] = 32'b00000011011010010010111011111000;
   assign mem[308575:308544] = 32'b11111110000000011001001100110110;
   assign mem[308607:308576] = 32'b11111101100101010100111010101000;
   assign mem[308639:308608] = 32'b00000011100100001011011110101100;
   assign mem[308671:308640] = 32'b00000100110000101001011111110000;
   assign mem[308703:308672] = 32'b11101111111001110111000101100000;
   assign mem[308735:308704] = 32'b00000010111101100111010100101000;
   assign mem[308767:308736] = 32'b00000111000011011100000111001000;
   assign mem[308799:308768] = 32'b11111010010101101111111000110000;
   assign mem[308831:308800] = 32'b00000100011000101100000001101000;
   assign mem[308863:308832] = 32'b11101101101010001001001010000000;
   assign mem[308895:308864] = 32'b00000110101101100001110011011000;
   assign mem[308927:308896] = 32'b11111000101110111011111111101000;
   assign mem[308959:308928] = 32'b11111111010011110000001111101011;
   assign mem[308991:308960] = 32'b00000000001110100101110101110111;
   assign mem[309023:308992] = 32'b11111011101010111100111111111000;
   assign mem[309055:309024] = 32'b11111101111111010000110010101100;
   assign mem[309087:309056] = 32'b00000001000101011101101100001110;
   assign mem[309119:309088] = 32'b00000010010110100111001100011100;
   assign mem[309151:309120] = 32'b00000100110000011011101011111000;
   assign mem[309183:309152] = 32'b00000001101100101111001101001110;
   assign mem[309215:309184] = 32'b00000110010000001101000100101000;
   assign mem[309247:309216] = 32'b11111011111000011101001110100000;
   assign mem[309279:309248] = 32'b11110111110011110110011111110000;
   assign mem[309311:309280] = 32'b11110011100010111001000011010000;
   assign mem[309343:309312] = 32'b11111111110111010100010101001101;
   assign mem[309375:309344] = 32'b00001000001100111001101010010000;
   assign mem[309407:309376] = 32'b11111011001000001100000101011000;
   assign mem[309439:309408] = 32'b00000101000101111000111010100000;
   assign mem[309471:309440] = 32'b00000001111011100101110011100010;
   assign mem[309503:309472] = 32'b00001001001001011100010010100000;
   assign mem[309535:309504] = 32'b11111011101111001010010001000000;
   assign mem[309567:309536] = 32'b11110111110011110010101001110000;
   assign mem[309599:309568] = 32'b00000010101110011011100101100100;
   assign mem[309631:309600] = 32'b00000011111101111110100010000100;
   assign mem[309663:309632] = 32'b11111101111111010011011100110100;
   assign mem[309695:309664] = 32'b00000110111110010100110111001000;
   assign mem[309727:309696] = 32'b11111111000100000011011110011101;
   assign mem[309759:309728] = 32'b11110111110100101011000110100000;
   assign mem[309791:309760] = 32'b11101010100101100010111000100000;
   assign mem[309823:309792] = 32'b00000111000001110101010010111000;
   assign mem[309855:309824] = 32'b11111111001011001101010010100100;
   assign mem[309887:309856] = 32'b00000111001100100010000001001000;
   assign mem[309919:309888] = 32'b11111111001011011001000010101110;
   assign mem[309951:309920] = 32'b00001000010101000100111010010000;
   assign mem[309983:309952] = 32'b11101110011110001000110000100000;
   assign mem[310015:309984] = 32'b11111011111010100000011100011000;
   assign mem[310047:310016] = 32'b00000011011111101110001101101000;
   assign mem[310079:310048] = 32'b11111111001111011100110000011011;
   assign mem[310111:310080] = 32'b00000100110110100111111111010000;
   assign mem[310143:310112] = 32'b11111101000001010011111110001100;
   assign mem[310175:310144] = 32'b00000001101010110000010101110100;
   assign mem[310207:310176] = 32'b11111001010101110101111111000000;
   assign mem[310239:310208] = 32'b11111110000011111000110001010000;
   assign mem[310271:310240] = 32'b00000010011011010000001010000000;
   assign mem[310303:310272] = 32'b00000010010110110001010010001000;
   assign mem[310335:310304] = 32'b11110111101111010001001001010000;
   assign mem[310367:310336] = 32'b00000010000000111011010000101000;
   assign mem[310399:310368] = 32'b11111111000110111110011001011010;
   assign mem[310431:310400] = 32'b11111100110000111001010110101100;
   assign mem[310463:310432] = 32'b00000000011110001101000000010010;
   assign mem[310495:310464] = 32'b00000011110100000110100111110100;
   assign mem[310527:310496] = 32'b11111101011000100110101110110100;
   assign mem[310559:310528] = 32'b00000001000011110010111010101110;
   assign mem[310591:310560] = 32'b00000110010011110100111001010000;
   assign mem[310623:310592] = 32'b11111011111100100111001100101000;
   assign mem[310655:310624] = 32'b00000000100100000010101100110011;
   assign mem[310687:310656] = 32'b11111011101111001111000001000000;
   assign mem[310719:310688] = 32'b11110000111000010010001101010000;
   assign mem[310751:310720] = 32'b00000101111001110000011001101000;
   assign mem[310783:310752] = 32'b11111011000000110110000011101000;
   assign mem[310815:310784] = 32'b11111011011101101101010011010000;
   assign mem[310847:310816] = 32'b11111101101110110101000010001100;
   assign mem[310879:310848] = 32'b00000001000101111101101110010100;
   assign mem[310911:310880] = 32'b11111111110000110100001111000100;
   assign mem[310943:310912] = 32'b00000110001011000010111011110000;
   assign mem[310975:310944] = 32'b11111011101010011110001100111000;
   assign mem[311007:310976] = 32'b00000011111110101101111011110100;
   assign mem[311039:311008] = 32'b11111111111110010111100100110100;
   assign mem[311071:311040] = 32'b11111010100000101100100011110000;
   assign mem[311103:311072] = 32'b00000111010111110001101000010000;
   assign mem[311135:311104] = 32'b11111111111000110110000010010010;
   assign mem[311167:311136] = 32'b00000010100001011111010010110100;
   assign mem[311199:311168] = 32'b11111011010100111010010011110000;
   assign mem[311231:311200] = 32'b11111110110101101010101011110110;
   assign mem[311263:311232] = 32'b11111110011101100010111000010000;
   assign mem[311295:311264] = 32'b11111111001011100010010100100100;
   assign mem[311327:311296] = 32'b11111000110101001000011101000000;
   assign mem[311359:311328] = 32'b00000001000001100000110000010000;
   assign mem[311391:311360] = 32'b11111011010010001101010100001000;
   assign mem[311423:311392] = 32'b00000100000011010111101101100000;
   assign mem[311455:311424] = 32'b11111110011001001100000100010010;
   assign mem[311487:311456] = 32'b00000111000011001000001000000000;
   assign mem[311519:311488] = 32'b11101110101101010010011010100000;
   assign mem[311551:311520] = 32'b00000011011000001001110111100000;
   assign mem[311583:311552] = 32'b11110011110001100101100110000000;
   assign mem[311615:311584] = 32'b11110111111101010011011100010000;
   assign mem[311647:311616] = 32'b11111011001010001010000011100000;
   assign mem[311679:311648] = 32'b00000010001111001101010000100000;
   assign mem[311711:311680] = 32'b00000111000111100111011110000000;
   assign mem[311743:311712] = 32'b11111111011101001010111100000110;
   assign mem[311775:311744] = 32'b00000011111101000000011110101100;
   assign mem[311807:311776] = 32'b11111111000001100110011011001111;
   assign mem[311839:311808] = 32'b00000111001101100001111100001000;
   assign mem[311871:311840] = 32'b11111100100100001100100111110000;
   assign mem[311903:311872] = 32'b11111110111110100000101011111110;
   assign mem[311935:311904] = 32'b11110011000100011111110100110000;
   assign mem[311967:311936] = 32'b11110110100000111101010001010000;
   assign mem[311999:311968] = 32'b11111100000110010110111100011100;
   assign mem[312031:312000] = 32'b00000110000101011110001001111000;
   assign mem[312063:312032] = 32'b11111001100100000011101111110000;
   assign mem[312095:312064] = 32'b00000000011011110011100010100000;
   assign mem[312127:312096] = 32'b11111010110010000010110110010000;
   assign mem[312159:312128] = 32'b11111110001011011011001101011100;
   assign mem[312191:312160] = 32'b11111010100111100010001010110000;
   assign mem[312223:312192] = 32'b00000011001010010001000000010100;
   assign mem[312255:312224] = 32'b11111101011111100111000001100100;
   assign mem[312287:312256] = 32'b00000110111111110110100110011000;
   assign mem[312319:312288] = 32'b11111011000010110101001010111000;
   assign mem[312351:312320] = 32'b11111011101000001100110101101000;
   assign mem[312383:312352] = 32'b00001000001010000101111000100000;
   assign mem[312415:312384] = 32'b00000010011000100000010011001100;
   assign mem[312447:312416] = 32'b11111110001110001010001000001000;
   assign mem[312479:312448] = 32'b00000110101010101100111000000000;
   assign mem[312511:312480] = 32'b00000000111110001101010110111011;
   assign mem[312543:312512] = 32'b11111100110111000011101001100100;
   assign mem[312575:312544] = 32'b11111110111011100001000001010110;
   assign mem[312607:312576] = 32'b11111000100001010111110011011000;
   assign mem[312639:312608] = 32'b11111010100100000110100000100000;
   assign mem[312671:312640] = 32'b00000000011000000100000111110010;
   assign mem[312703:312672] = 32'b11110110010001100011100010010000;
   assign mem[312735:312704] = 32'b00000000100100101100100101010010;
   assign mem[312767:312736] = 32'b00000010001101110101110011001100;
   assign mem[312799:312768] = 32'b00000001110110011011111001111100;
   assign mem[312831:312800] = 32'b11111011101110101100110000101000;
   assign mem[312863:312832] = 32'b00000100100101111100110101011000;
   assign mem[312895:312864] = 32'b11111101010111100111001111101100;
   assign mem[312927:312896] = 32'b11111100110101111101111001010000;
   assign mem[312959:312928] = 32'b11111011101011100000000000001000;
   assign mem[312991:312960] = 32'b11111001010001001100010110100000;
   assign mem[313023:312992] = 32'b11110111110010010011101011000000;
   assign mem[313055:313024] = 32'b11110110110110110101000000000000;
   assign mem[313087:313056] = 32'b00000001011101011101101100001010;
   assign mem[313119:313088] = 32'b00001111001001111010100111000000;
   assign mem[313151:313120] = 32'b00000011011110110100101100111100;
   assign mem[313183:313152] = 32'b11110000111111011011111011100000;
   assign mem[313215:313184] = 32'b00000101100011100011110010101000;
   assign mem[313247:313216] = 32'b00000100100010001110000100001000;
   assign mem[313279:313248] = 32'b11111110001110110101111011000100;
   assign mem[313311:313280] = 32'b11111110101000110000110100000110;
   assign mem[313343:313312] = 32'b00000110100010111101111001101000;
   assign mem[313375:313344] = 32'b00001100000000000011010010100000;
   assign mem[313407:313376] = 32'b11111101100010111110010001111000;
   assign mem[313439:313408] = 32'b11110101011100001110100111100000;
   assign mem[313471:313440] = 32'b11111101010101001110100011111100;
   assign mem[313503:313472] = 32'b11111110010011000100011111101000;
   assign mem[313535:313504] = 32'b00001011100110011011010101110000;
   assign mem[313567:313536] = 32'b00000001000110100010000010111110;
   assign mem[313599:313568] = 32'b11100111000000010111010010100000;
   assign mem[313631:313600] = 32'b00000011011100101110110101111000;
   assign mem[313663:313632] = 32'b11110110011000011001110000110000;
   assign mem[313695:313664] = 32'b00000001010101110111110000001110;
   assign mem[313727:313696] = 32'b11111001011101110000111001101000;
   assign mem[313759:313728] = 32'b00000011111110000110011110010100;
   assign mem[313791:313760] = 32'b11110011101100110101111010110000;
   assign mem[313823:313792] = 32'b00000100010101100001100001001000;
   assign mem[313855:313824] = 32'b00000100010110000111000101111000;
   assign mem[313887:313856] = 32'b11111110011010001001100000001010;
   assign mem[313919:313888] = 32'b00000111111101100011010111101000;
   assign mem[313951:313920] = 32'b11110010011010101110111010010000;
   assign mem[313983:313952] = 32'b00000010110001010000110001101000;
   assign mem[314015:313984] = 32'b00000101101011100110111100000000;
   assign mem[314047:314016] = 32'b11111000111011101110101101010000;
   assign mem[314079:314048] = 32'b11111100011010001001100100000000;
   assign mem[314111:314080] = 32'b11111011001000010111011101010000;
   assign mem[314143:314112] = 32'b11111001100111010001100111000000;
   assign mem[314175:314144] = 32'b00000001010011100010110101111110;
   assign mem[314207:314176] = 32'b00000100000010010101000110000000;
   assign mem[314239:314208] = 32'b11111010001001111001100101000000;
   assign mem[314271:314240] = 32'b00001010011101010110010110010000;
   assign mem[314303:314272] = 32'b11111101010110101110101100101000;
   assign mem[314335:314304] = 32'b11111111111100011010000011010011;
   assign mem[314367:314336] = 32'b11110010101010111000010011100000;
   assign mem[314399:314368] = 32'b00000101011111000111000101101000;
   assign mem[314431:314400] = 32'b11111111110010010000100011000111;
   assign mem[314463:314432] = 32'b00000000100111101010001001011111;
   assign mem[314495:314464] = 32'b00000111111001011000111000111000;
   assign mem[314527:314496] = 32'b11111111101000110110011010111111;
   assign mem[314559:314528] = 32'b11111001100000000010100101110000;
   assign mem[314591:314560] = 32'b00000010110000101100111010010000;
   assign mem[314623:314592] = 32'b11110011000000111010001011110000;
   assign mem[314655:314624] = 32'b11111110111001000000111010000000;
   assign mem[314687:314656] = 32'b00000101000111100000011011111000;
   assign mem[314719:314688] = 32'b00000001010001010111001111001100;
   assign mem[314751:314720] = 32'b11111111000111000100110010110110;
   assign mem[314783:314752] = 32'b00000110001111111111101100011000;
   assign mem[314815:314784] = 32'b11111010101010011111100001111000;
   assign mem[314847:314816] = 32'b11111100110000011101110110010100;
   assign mem[314879:314848] = 32'b11111101101011011110100100001000;
   assign mem[314911:314880] = 32'b00000100101000001011001001111000;
   assign mem[314943:314912] = 32'b11110000111001111011001010010000;
   assign mem[314975:314944] = 32'b11111010111100011110000111000000;
   assign mem[315007:314976] = 32'b00000101101010001011010100011000;
   assign mem[315039:315008] = 32'b11111101011111100101000010000000;
   assign mem[315071:315040] = 32'b00000011100001100111101011000100;
   assign mem[315103:315072] = 32'b00000101100000010101111001000000;
   assign mem[315135:315104] = 32'b11111011100011010111000100010000;
   assign mem[315167:315136] = 32'b11111101000100011010011001010000;
   assign mem[315199:315168] = 32'b00000000011000100110000001110010;
   assign mem[315231:315200] = 32'b00000001111000100010011001111000;
   assign mem[315263:315232] = 32'b00001011010010011011001110010000;
   assign mem[315295:315264] = 32'b11111000111011010100101101010000;
   assign mem[315327:315296] = 32'b00000011000100100000011010111000;
   assign mem[315359:315328] = 32'b11111101110001010010000101111000;
   assign mem[315391:315360] = 32'b11110001101110011110100010000000;
   assign mem[315423:315392] = 32'b11111001101010000111111001011000;
   assign mem[315455:315424] = 32'b00001011011000111111111011000000;
   assign mem[315487:315456] = 32'b11110110011010010011001010110000;
   assign mem[315519:315488] = 32'b11111100000011110010100001110100;
   assign mem[315551:315520] = 32'b00000101110111100100001110010000;
   assign mem[315583:315552] = 32'b11101011111001101000110011100000;
   assign mem[315615:315584] = 32'b11110110111110111101000000110000;
   assign mem[315647:315616] = 32'b00000000100000101010110000101110;
   assign mem[315679:315648] = 32'b11111000111110101011111111000000;
   assign mem[315711:315680] = 32'b11110000101000111001000110000000;
   assign mem[315743:315712] = 32'b00000001011001110110110011101010;
   assign mem[315775:315744] = 32'b11111110000101011001111110110000;
   assign mem[315807:315776] = 32'b11111011011101000010101001110000;
   assign mem[315839:315808] = 32'b00001000101010100000010111100000;
   assign mem[315871:315840] = 32'b11111011101101011110011001001000;
   assign mem[315903:315872] = 32'b00000001010100000010110001101110;
   assign mem[315935:315904] = 32'b00000100100100110101000111110000;
   assign mem[315967:315936] = 32'b11111001101010001001000111010000;
   assign mem[315999:315968] = 32'b11111101000011101110110101001000;
   assign mem[316031:316000] = 32'b11111111001011110100101010011001;
   assign mem[316063:316032] = 32'b11111101101110011010010000010000;
   assign mem[316095:316064] = 32'b11111110100001111110010010110010;
   assign mem[316127:316096] = 32'b00000101111100000111101000100000;
   assign mem[316159:316128] = 32'b11110111000101100011100110100000;
   assign mem[316191:316160] = 32'b11111100010100100111101101010100;
   assign mem[316223:316192] = 32'b11111111101011000100010100000001;
   assign mem[316255:316224] = 32'b00001100111100010101110111100000;
   assign mem[316287:316256] = 32'b11111100000110000000110011111100;
   assign mem[316319:316288] = 32'b00000001111001001011100001101100;
   assign mem[316351:316320] = 32'b11111101100001000010000110011000;
   assign mem[316383:316352] = 32'b11111110000101001101011001111010;
   assign mem[316415:316384] = 32'b11110100111100001000110000010000;
   assign mem[316447:316416] = 32'b11111010001001001111000100011000;
   assign mem[316479:316448] = 32'b11111111011010010001010100100010;
   assign mem[316511:316480] = 32'b11101101000001011000101010000000;
   assign mem[316543:316512] = 32'b00000110101100101111011001011000;
   assign mem[316575:316544] = 32'b00000100111110011111000100111000;
   assign mem[316607:316576] = 32'b00000011101011110011101100010100;
   assign mem[316639:316608] = 32'b11110100100010000110010100100000;
   assign mem[316671:316640] = 32'b00000111011111000010101000111000;
   assign mem[316703:316672] = 32'b11110101100100001100100001000000;
   assign mem[316735:316704] = 32'b11111111011111001101100000010010;
   assign mem[316767:316736] = 32'b11111100101010100001101101110100;
   assign mem[316799:316768] = 32'b11111010110110111111100000001000;
   assign mem[316831:316800] = 32'b00000001011110101110000010100000;
   assign mem[316863:316832] = 32'b11101101111110110010010100100000;
   assign mem[316895:316864] = 32'b11111101110101100010000000010100;
   assign mem[316927:316896] = 32'b11111101001111101100110111001100;
   assign mem[316959:316928] = 32'b11111101001100110111010000011000;
   assign mem[316991:316960] = 32'b11111101111111010100000111011100;
   assign mem[317023:316992] = 32'b00000101010110000111000101011000;
   assign mem[317055:317024] = 32'b00001001011001010011001010000000;
   assign mem[317087:317056] = 32'b11111100100010001111000001111100;
   assign mem[317119:317088] = 32'b00000010000111001110100011000000;
   assign mem[317151:317120] = 32'b11111111011011000000001111100111;
   assign mem[317183:317152] = 32'b00000100100010110111101001111000;
   assign mem[317215:317184] = 32'b11111101010101011000100000000000;
   assign mem[317247:317216] = 32'b11111011010000101010001100110000;
   assign mem[317279:317248] = 32'b00000001011101010101110011111100;
   assign mem[317311:317280] = 32'b00000100111101001101110000001000;
   assign mem[317343:317312] = 32'b00000001001010110001000001010010;
   assign mem[317375:317344] = 32'b11111011010111110101110010000000;
   assign mem[317407:317376] = 32'b00000000111011010101001110010100;
   assign mem[317439:317408] = 32'b11111110110100110101011111111000;
   assign mem[317471:317440] = 32'b00001000001100100001010010110000;
   assign mem[317503:317472] = 32'b11110101101000001110011011100000;
   assign mem[317535:317504] = 32'b00000111011110000111111001100000;
   assign mem[317567:317536] = 32'b11110011000011000101000001110000;
   assign mem[317599:317568] = 32'b00000011110110011011011001111000;
   assign mem[317631:317600] = 32'b00000000000011011001001110000011;
   assign mem[317663:317632] = 32'b00000001101001110110111010110000;
   assign mem[317695:317664] = 32'b11110111111000001110010110110000;
   assign mem[317727:317696] = 32'b00000111110111010011010101001000;
   assign mem[317759:317728] = 32'b11110011000111110100111001010000;
   assign mem[317791:317760] = 32'b00000100111010111111111000101000;
   assign mem[317823:317792] = 32'b11101011010100000010100110100000;
   assign mem[317855:317824] = 32'b11111111100011000111010100101001;
   assign mem[317887:317856] = 32'b11110000100010010110001001100000;
   assign mem[317919:317888] = 32'b00000100010100111100111010100000;
   assign mem[317951:317920] = 32'b11111111000011011100001101001101;
   assign mem[317983:317952] = 32'b00000000011100111000111011001100;
   assign mem[318015:317984] = 32'b11111000011101010111101011100000;
   assign mem[318047:318016] = 32'b00000000011110010101101110111100;
   assign mem[318079:318048] = 32'b00001000000100000110101011010000;
   assign mem[318111:318080] = 32'b00000100101101010010100010010000;
   assign mem[318143:318112] = 32'b00000110100010010100001011100000;
   assign mem[318175:318144] = 32'b11111101110010110011001011111000;
   assign mem[318207:318176] = 32'b11111011111100000000010001010000;
   assign mem[318239:318208] = 32'b00000111001010111101101010011000;
   assign mem[318271:318240] = 32'b11110111110101000110110101000000;
   assign mem[318303:318272] = 32'b00000001011100000110111011110010;
   assign mem[318335:318304] = 32'b00000001100100101001001001001010;
   assign mem[318367:318336] = 32'b00000110110010000111100110100000;
   assign mem[318399:318368] = 32'b00000000110000011000000000011111;
   assign mem[318431:318400] = 32'b11110001010010011001011110100000;
   assign mem[318463:318432] = 32'b00000110100110000101110010000000;
   assign mem[318495:318464] = 32'b00000110100111000000000000010000;
   assign mem[318527:318496] = 32'b11111100001001110100000001001000;
   assign mem[318559:318528] = 32'b11111011110011001101111000001000;
   assign mem[318591:318560] = 32'b00000000111110110101010111100111;
   assign mem[318623:318592] = 32'b11111000110100011101100000100000;
   assign mem[318655:318624] = 32'b00000001110011000110101010001000;
   assign mem[318687:318656] = 32'b00001000010100110000101111100000;
   assign mem[318719:318688] = 32'b11110110111101111000001110000000;
   assign mem[318751:318720] = 32'b11111001010011010101011010100000;
   assign mem[318783:318752] = 32'b00000101111111110110111011011000;
   assign mem[318815:318784] = 32'b11110110001100101001100000010000;
   assign mem[318847:318816] = 32'b00000010110100011010001110000000;
   assign mem[318879:318848] = 32'b00000010011011110111110011010100;
   assign mem[318911:318880] = 32'b00000110011010110011110111111000;
   assign mem[318943:318912] = 32'b11101000001111001010100100100000;
   assign mem[318975:318944] = 32'b11111101111110100110010100011000;
   assign mem[319007:318976] = 32'b00000001011100001001011100101100;
   assign mem[319039:319008] = 32'b11111010011111100111011010111000;
   assign mem[319071:319040] = 32'b11111011010101001101111101101000;
   assign mem[319103:319072] = 32'b11111000111101000010001100110000;
   assign mem[319135:319104] = 32'b00000010010111111110000001101000;
   assign mem[319167:319136] = 32'b00000111000001010001011100011000;
   assign mem[319199:319168] = 32'b11110011100011101110100011010000;
   assign mem[319231:319200] = 32'b00001010000001100011010010100000;
   assign mem[319263:319232] = 32'b11110010001100001010101001110000;
   assign mem[319295:319264] = 32'b11110101000001110110011110010000;
   assign mem[319327:319296] = 32'b11111010110001000110001001101000;
   assign mem[319359:319328] = 32'b11111011001101011001000011001000;
   assign mem[319391:319360] = 32'b11111101011101010111101001000100;
   assign mem[319423:319392] = 32'b11111100110110000110001110010100;
   assign mem[319455:319424] = 32'b00000110110101011010101000000000;
   assign mem[319487:319456] = 32'b00000000101100101111001111011100;
   assign mem[319519:319488] = 32'b00000101110000111010101000100000;
   assign mem[319551:319520] = 32'b11111001111011101001110110010000;
   assign mem[319583:319552] = 32'b00000000111001100011000010100110;
   assign mem[319615:319584] = 32'b11110100111011001101010111110000;
   assign mem[319647:319616] = 32'b11111001101101010110100100010000;
   assign mem[319679:319648] = 32'b00000010010110111110011111101100;
   assign mem[319711:319680] = 32'b11101110011000011001010001100000;
   assign mem[319743:319712] = 32'b00000111010011110001110110101000;
   assign mem[319775:319744] = 32'b11111111101100010101101010010100;
   assign mem[319807:319776] = 32'b00000001001101000001111011101000;
   assign mem[319839:319808] = 32'b00000001001100101111001101111010;
   assign mem[319871:319840] = 32'b00000010011100111010101000101000;
   assign mem[319903:319872] = 32'b11101100010101110010010110000000;
   assign mem[319935:319904] = 32'b00000101100011011111001111101000;
   assign mem[319967:319936] = 32'b11111111000000110111000001001001;
   assign mem[319999:319968] = 32'b11111011111010101010110000010000;
   assign mem[320031:320000] = 32'b00000011010011011101010010010100;
   assign mem[320063:320032] = 32'b11101101101000000010100010100000;
   assign mem[320095:320064] = 32'b11111011110010100101100001000000;
   assign mem[320127:320096] = 32'b11110111101110010110001000110000;
   assign mem[320159:320128] = 32'b00000101101110000101100100101000;
   assign mem[320191:320160] = 32'b11111011101101010011010110000000;
   assign mem[320223:320192] = 32'b00000100110010000110100101010000;
   assign mem[320255:320224] = 32'b11111000100110110011110110000000;
   assign mem[320287:320256] = 32'b00000011100011111000000001101000;
   assign mem[320319:320288] = 32'b00000100101100010011011011100000;
   assign mem[320351:320320] = 32'b11111101010110010101100011010000;
   assign mem[320383:320352] = 32'b00000100010101010111110000011000;
   assign mem[320415:320384] = 32'b11111001101101100111011010111000;
   assign mem[320447:320416] = 32'b11111110100100100110001110010100;
   assign mem[320479:320448] = 32'b00000010101111010110011101011100;
   assign mem[320511:320480] = 32'b00000101010011010000001110100000;
   assign mem[320543:320512] = 32'b11110011100111000010011000110000;
   assign mem[320575:320544] = 32'b00000100101001100110110110110000;
   assign mem[320607:320576] = 32'b11111011011100001011001101011000;
   assign mem[320639:320608] = 32'b11111011101001111111100100110000;
   assign mem[320671:320640] = 32'b11111100010111010001110010000100;
   assign mem[320703:320672] = 32'b00000000010100011001110101000010;
   assign mem[320735:320704] = 32'b11111100000000000000011110010100;
   assign mem[320767:320736] = 32'b11111101000111101110100101011100;
   assign mem[320799:320768] = 32'b00000010110001111011000010100100;
   assign mem[320831:320800] = 32'b11111101101101110111100101110100;
   assign mem[320863:320832] = 32'b11111110101000010110101010110000;
   assign mem[320895:320864] = 32'b11111110000011010100110000000000;
   assign mem[320927:320896] = 32'b00000000010111001110000000000111;
   assign mem[320959:320928] = 32'b00000010011110101001010010001100;
   assign mem[320991:320960] = 32'b11111011111111000001111101110000;
   assign mem[321023:320992] = 32'b11111110101111110001001011100100;
   assign mem[321055:321024] = 32'b00000010111001101000111101111100;
   assign mem[321087:321056] = 32'b00000111101010000100010111100000;
   assign mem[321119:321088] = 32'b00000100011001111110001100101000;
   assign mem[321151:321120] = 32'b11111000000111101101111000101000;
   assign mem[321183:321152] = 32'b11111011111111011111111110110000;
   assign mem[321215:321184] = 32'b11110101101011111000000001010000;
   assign mem[321247:321216] = 32'b11111110101110011110011100100100;
   assign mem[321279:321248] = 32'b00000100010111101010000111001000;
   assign mem[321311:321280] = 32'b00000100011111001101111110100000;
   assign mem[321343:321312] = 32'b11111000100001111011101000100000;
   assign mem[321375:321344] = 32'b00000110111111110010010100110000;
   assign mem[321407:321376] = 32'b11111100110100101011001111010100;
   assign mem[321439:321408] = 32'b11111110001010101010100101101000;
   assign mem[321471:321440] = 32'b11110011111001011000101101010000;
   assign mem[321503:321472] = 32'b00000100001110001101111100111000;
   assign mem[321535:321504] = 32'b11110101001110001010100010100000;
   assign mem[321567:321536] = 32'b00000111001011000100100101011000;
   assign mem[321599:321568] = 32'b00000001101101100000010001010110;
   assign mem[321631:321600] = 32'b00000011001100001001110110010100;
   assign mem[321663:321632] = 32'b11111101110011110111000010001100;
   assign mem[321695:321664] = 32'b00000100001101110110110111010000;
   assign mem[321727:321696] = 32'b00000011001010101101010011010000;
   assign mem[321759:321728] = 32'b11111100001111100110100010000000;
   assign mem[321791:321760] = 32'b00000010110001110000110110110000;
   assign mem[321823:321792] = 32'b11111011000010100101100110101000;
   assign mem[321855:321824] = 32'b11111011100100001110001110010000;
   assign mem[321887:321856] = 32'b00000101100111111010010000111000;
   assign mem[321919:321888] = 32'b11111011101000000110111000111000;
   assign mem[321951:321920] = 32'b00000100110001010011101001101000;
   assign mem[321983:321952] = 32'b11111000000000010010001101000000;
   assign mem[322015:321984] = 32'b00000010010011001001101100010100;
   assign mem[322047:322016] = 32'b11110111110110100000000000110000;
   assign mem[322079:322048] = 32'b11111100100110000101010011101100;
   assign mem[322111:322080] = 32'b11111011111110011000101110101000;
   assign mem[322143:322112] = 32'b00001001000110100101011001110000;
   assign mem[322175:322144] = 32'b11110010110101101100101101010000;
   assign mem[322207:322176] = 32'b00000000010010000101110001001011;
   assign mem[322239:322208] = 32'b00000011111100111110011100110100;
   assign mem[322271:322240] = 32'b11111111000101000101110001011010;
   assign mem[322303:322272] = 32'b11111101111101010100000010111000;
   assign mem[322335:322304] = 32'b00000000000111000001010000011000;
   assign mem[322367:322336] = 32'b11111100111001011001101001100100;
   assign mem[322399:322368] = 32'b11111100000111001110111100111100;
   assign mem[322431:322400] = 32'b11111101110100000001000100100000;
   assign mem[322463:322432] = 32'b00000001011010101010111000010010;
   assign mem[322495:322464] = 32'b00000001000111000100011011100110;
   assign mem[322527:322496] = 32'b00000011000101001001001010001100;
   assign mem[322559:322528] = 32'b00000010010101000000001101110100;
   assign mem[322591:322560] = 32'b00000001101011000101001011000010;
   assign mem[322623:322592] = 32'b11110111110101000001110101000000;
   assign mem[322655:322624] = 32'b11111110000011111101011101010010;
   assign mem[322687:322656] = 32'b11111101010110110100011111100000;
   assign mem[322719:322688] = 32'b00000011100100101010110000001000;
   assign mem[322751:322720] = 32'b11111100110111100101000111110100;
   assign mem[322783:322752] = 32'b00000000011101010101111100000000;
   assign mem[322815:322784] = 32'b11111101010001100000110110010000;
   assign mem[322847:322816] = 32'b11111110101111110000011011101100;
   assign mem[322879:322848] = 32'b11111101111111000111001111001000;
   assign mem[322911:322880] = 32'b00000011110111111011010100101100;
   assign mem[322943:322912] = 32'b11111011110111000100111110011000;
   assign mem[322975:322944] = 32'b00000010101101100101111111011000;
   assign mem[323007:322976] = 32'b11110110111010010110100000010000;
   assign mem[323039:323008] = 32'b00000001111000000001110011000100;
   assign mem[323071:323040] = 32'b11111010111111110010010111000000;
   assign mem[323103:323072] = 32'b00000100011010001110010110100000;
   assign mem[323135:323104] = 32'b11111010111111101110010000101000;
   assign mem[323167:323136] = 32'b00000010000010000100100111101000;
   assign mem[323199:323168] = 32'b11110110110101110011010010100000;
   assign mem[323231:323200] = 32'b00001001111111111001010001010000;
   assign mem[323263:323232] = 32'b11111110011011110000001111010000;
   assign mem[323295:323264] = 32'b00000001101010111111010100000100;
   assign mem[323327:323296] = 32'b11101111011010011101001101100000;
   assign mem[323359:323328] = 32'b00000111111010100100111000101000;
   assign mem[323391:323360] = 32'b00000001101100101101100000110110;
   assign mem[323423:323392] = 32'b11111111101000111000010000110101;
   assign mem[323455:323424] = 32'b11111011010110001110100011001000;
   assign mem[323487:323456] = 32'b00000110110010110101100011100000;
   assign mem[323519:323488] = 32'b11111011001101110010000001111000;
   assign mem[323551:323520] = 32'b00000001010100110111010011010110;
   assign mem[323583:323552] = 32'b11111110010100111100001101000010;
   assign mem[323615:323584] = 32'b11111101010010111101110100010100;
   assign mem[323647:323616] = 32'b11111111101111100110000010100100;
   assign mem[323679:323648] = 32'b11111101100110101110010000111000;
   assign mem[323711:323680] = 32'b00000001010100001011101001110100;
   assign mem[323743:323712] = 32'b00000001101000001100111111000000;
   assign mem[323775:323744] = 32'b00000010011110111000001101110000;
   assign mem[323807:323776] = 32'b00000010110101001010000010011100;
   assign mem[323839:323808] = 32'b00000010000111100001110111110100;
   assign mem[323871:323840] = 32'b00000100010111001010110101101000;
   assign mem[323903:323872] = 32'b00000111000111110001101000011000;
   assign mem[323935:323904] = 32'b11111110001100001001100011001000;
   assign mem[323967:323936] = 32'b11111001001001111111111011001000;
   assign mem[323999:323968] = 32'b00000101101001001000110011100000;
   assign mem[324031:324000] = 32'b11111100100010001111010000000100;
   assign mem[324063:324032] = 32'b11111000101011101000100101110000;
   assign mem[324095:324064] = 32'b11111100111001011110010111011000;
   assign mem[324127:324096] = 32'b11111101011111101111111010101100;
   assign mem[324159:324128] = 32'b00000001100101001111100010110100;
   assign mem[324191:324160] = 32'b00000010011011010010010010100000;
   assign mem[324223:324192] = 32'b00000011111011000000001110100100;
   assign mem[324255:324224] = 32'b11111101011100000001011011000100;
   assign mem[324287:324256] = 32'b11111111000001000111010001110111;
   assign mem[324319:324288] = 32'b11111110101111011101011101000010;
   assign mem[324351:324320] = 32'b11111111110101110110001011001101;
   assign mem[324383:324352] = 32'b11111010011011010001101011111000;
   assign mem[324415:324384] = 32'b11111010000011000110100011001000;
   assign mem[324447:324416] = 32'b11111011100010101000110011100000;
   assign mem[324479:324448] = 32'b00000100100101000001000111011000;
   assign mem[324511:324480] = 32'b00000010010010101001000000100100;
   assign mem[324543:324512] = 32'b11111001110110110100011011001000;
   assign mem[324575:324544] = 32'b00000100101100000010110010110000;
   assign mem[324607:324576] = 32'b11110111100110010000000000100000;
   assign mem[324639:324608] = 32'b00000100111100000111100000110000;
   assign mem[324671:324640] = 32'b00000011111010011001010110011000;
   assign mem[324703:324672] = 32'b11111100010011001010101011011100;
   assign mem[324735:324704] = 32'b00000000010111111001011110001101;
   assign mem[324767:324736] = 32'b00000001101010010001010101110010;
   assign mem[324799:324768] = 32'b11111110100011001010001101001110;
   assign mem[324831:324800] = 32'b11111110100000100001010101101110;
   assign mem[324863:324832] = 32'b11111010101100110100011100001000;
   assign mem[324895:324864] = 32'b00001001100001011101010101110000;
   assign mem[324927:324896] = 32'b11111111001100111100101110001000;
   assign mem[324959:324928] = 32'b00000001100001100111100001010100;
   assign mem[324991:324960] = 32'b11111110001101010110011010101010;
   assign mem[325023:324992] = 32'b11111110010000011100000001010100;
   assign mem[325055:325024] = 32'b11111100110111010010101110100100;
   assign mem[325087:325056] = 32'b00000011101011011101011111101000;
   assign mem[325119:325088] = 32'b00000000000101110000010010010111;
   assign mem[325151:325120] = 32'b00000010101010001011001000010100;
   assign mem[325183:325152] = 32'b11111110110010001100010101001000;
   assign mem[325215:325184] = 32'b00000110101101001111110010111000;
   assign mem[325247:325216] = 32'b11111110100011110001011111111100;
   assign mem[325279:325248] = 32'b11111111001100011000111010110111;
   assign mem[325311:325280] = 32'b11111011011010000011111011100000;
   assign mem[325343:325312] = 32'b11111110011000010110000100010110;
   assign mem[325375:325344] = 32'b11111010110111100111001111111000;
   assign mem[325407:325376] = 32'b00000000111010001111110010111111;
   assign mem[325439:325408] = 32'b11111110010001111001110110111000;
   assign mem[325471:325440] = 32'b00000100011000001000010011101000;
   assign mem[325503:325472] = 32'b11111011101001110011011001000000;
   assign mem[325535:325504] = 32'b11111000101100101010011100011000;
   assign mem[325567:325536] = 32'b11111010101100001111111001111000;
   assign mem[325599:325568] = 32'b00000111010111101000011001100000;
   assign mem[325631:325600] = 32'b11111101011101001001101100001000;
   assign mem[325663:325632] = 32'b00000101111111101101010100110000;
   assign mem[325695:325664] = 32'b11110100101100011001110100110000;
   assign mem[325727:325696] = 32'b00000011011100000111001011111000;
   assign mem[325759:325728] = 32'b00000110001001111110111100010000;
   assign mem[325791:325760] = 32'b11111000011011110001000111101000;
   assign mem[325823:325792] = 32'b00000110100100111001110110100000;
   assign mem[325855:325824] = 32'b11111100011000011111000001000000;
   assign mem[325887:325856] = 32'b00000111101011111100011111100000;
   assign mem[325919:325888] = 32'b11111010110010011010110010101000;
   assign mem[325951:325920] = 32'b00000101001011000110011111110000;
   assign mem[325983:325952] = 32'b11110001011010111101101011110000;
   assign mem[326015:325984] = 32'b11110111010111011111101100110000;
   assign mem[326047:326016] = 32'b00000000001001110100100010101110;
   assign mem[326079:326048] = 32'b11110100101110110010110111010000;
   assign mem[326111:326080] = 32'b00000000100101010000001011101011;
   assign mem[326143:326112] = 32'b11111011100100010011110101101000;
   assign mem[326175:326144] = 32'b00000100101011110101110110011000;
   assign mem[326207:326176] = 32'b00000110101011100011111100000000;
   assign mem[326239:326208] = 32'b11110110100110110110010100010000;
   assign mem[326271:326240] = 32'b00000001101011110010101000010100;
   assign mem[326303:326272] = 32'b11110110101011101001110111000000;
   assign mem[326335:326304] = 32'b11111010000100110001110011100000;
   assign mem[326367:326336] = 32'b00000101111001100110001000010000;
   assign mem[326399:326368] = 32'b11101100111010101100101100100000;
   assign mem[326431:326400] = 32'b11101111100101100001011111100000;
   assign mem[326463:326432] = 32'b00000100101110110100001001000000;
   assign mem[326495:326464] = 32'b00000011001001001001100000100000;
   assign mem[326527:326496] = 32'b00000001001000110011000000110100;
   assign mem[326559:326528] = 32'b00000001010111110000100101010110;
   assign mem[326591:326560] = 32'b11111111010100110111010100011001;
   assign mem[326623:326592] = 32'b11110111110101101000110011110000;
   assign mem[326655:326624] = 32'b00000000111001010100001000001011;
   assign mem[326687:326656] = 32'b00000010101011110011101011110100;
   assign mem[326719:326688] = 32'b11110001000000000001001000100000;
   assign mem[326751:326720] = 32'b00000110100110011001011000111000;
   assign mem[326783:326752] = 32'b11110010111111110110101010000000;
   assign mem[326815:326784] = 32'b00000100111100100101100001000000;
   assign mem[326847:326816] = 32'b11110000110111011101010000000000;
   assign mem[326879:326848] = 32'b00000001100001110001100101111010;
   assign mem[326911:326880] = 32'b11111011010111111111001000100000;
   assign mem[326943:326912] = 32'b11111111101010010111100011000011;
   assign mem[326975:326944] = 32'b11111101001010010000111101010100;
   assign mem[327007:326976] = 32'b00000100011101111100110000001000;
   assign mem[327039:327008] = 32'b11111100000101001111100011111100;
   assign mem[327071:327040] = 32'b00000010001001111011001001001100;
   assign mem[327103:327072] = 32'b11111001111110010010110100100000;
   assign mem[327135:327104] = 32'b00000011001100110100001000110100;
   assign mem[327167:327136] = 32'b00000001110110010110010011111000;
   assign mem[327199:327168] = 32'b11111001010111100111010001101000;
   assign mem[327231:327200] = 32'b11111100000101100011010001010100;
   assign mem[327263:327232] = 32'b00000010101000101011101111110100;
   assign mem[327295:327264] = 32'b11111011001001011100011111111000;
   assign mem[327327:327296] = 32'b11111111101101100001000111111110;
   assign mem[327359:327328] = 32'b00000000100011111011011110101011;
   assign mem[327391:327360] = 32'b00000011100110100010110000011100;
   assign mem[327423:327392] = 32'b11111011110111001100101010111000;
   assign mem[327455:327424] = 32'b00000001111010011110011111110000;
   assign mem[327487:327456] = 32'b11110101011110111000110001000000;
   assign mem[327519:327488] = 32'b11111001110100000111111100000000;
   assign mem[327551:327520] = 32'b11111110001001111100000001111010;
   assign mem[327583:327552] = 32'b00000100000101001110100000101000;
   assign mem[327615:327584] = 32'b11111010010110100110100011000000;
   assign mem[327647:327616] = 32'b00000001001010001011110000100100;
   assign mem[327679:327648] = 32'b00000001111110010011011111011100;
   assign mem[327711:327680] = 32'b11111011010000101010011111010000;
   assign mem[327743:327712] = 32'b11111110010010001011000000011000;
   assign mem[327775:327744] = 32'b11111100001001001111011000011100;
   assign mem[327807:327776] = 32'b00000000010010000110100110110001;
   assign mem[327839:327808] = 32'b00000001100000110001101111100100;
   assign mem[327871:327840] = 32'b00000001111000000001110001001110;
   assign mem[327903:327872] = 32'b11111110001101011001110010001100;
   assign mem[327935:327904] = 32'b11111101000001001100001011001000;
   assign mem[327967:327936] = 32'b11111111101111011110010010000011;
   assign mem[327999:327968] = 32'b00000011010010000001111100100100;
   assign mem[328031:328000] = 32'b00000000011111100110110101100100;
   assign mem[328063:328032] = 32'b00000010011011111110111001011000;
   assign mem[328095:328064] = 32'b11100010110000100011011010000000;
   assign mem[328127:328096] = 32'b00001001010101110011111011110000;
   assign mem[328159:328128] = 32'b11111001011000001110110010010000;
   assign mem[328191:328160] = 32'b00000111111010100101010011110000;
   assign mem[328223:328192] = 32'b11101100000000000001111111000000;
   assign mem[328255:328224] = 32'b00001011101010110100110011100000;
   assign mem[328287:328256] = 32'b11100110001110110000001110000000;
   assign mem[328319:328288] = 32'b00000001001001010111011010111110;
   assign mem[328351:328320] = 32'b00000010001110001011101110011000;
   assign mem[328383:328352] = 32'b11110111101101101001101110000000;
   assign mem[328415:328384] = 32'b11111100111010000001001010001100;
   assign mem[328447:328416] = 32'b11111010100000100100001000100000;
   assign mem[328479:328448] = 32'b00000100000110010001110101010000;
   assign mem[328511:328480] = 32'b00000010000100101000010110111100;
   assign mem[328543:328512] = 32'b00000000101101111010011000010010;
   assign mem[328575:328544] = 32'b11110001111000010011110101010000;
   assign mem[328607:328576] = 32'b00000111010101010111101101000000;
   assign mem[328639:328608] = 32'b11111111001110110010001100001000;
   assign mem[328671:328640] = 32'b11110101010101111011101100010000;
   assign mem[328703:328672] = 32'b11110110111110000111101100110000;
   assign mem[328735:328704] = 32'b11110100011011000010001100100000;
   assign mem[328767:328736] = 32'b00000011011010010011110010000000;
   assign mem[328799:328768] = 32'b00000101110011011010110000100000;
   assign mem[328831:328800] = 32'b11111110100000010010001001101000;
   assign mem[328863:328832] = 32'b11101010000100001011111011000000;
   assign mem[328895:328864] = 32'b11111110111101011111101010011010;
   assign mem[328927:328896] = 32'b11111011000011111101111110010000;
   assign mem[328959:328928] = 32'b00000110011000001011000001010000;
   assign mem[328991:328960] = 32'b11101100001001110110111000100000;
   assign mem[329023:328992] = 32'b00000011110000010111111110111000;
   assign mem[329055:329024] = 32'b11111111001001011110000101101111;
   assign mem[329087:329056] = 32'b00000011011011111011110111110000;
   assign mem[329119:329088] = 32'b00000011101110111110110001100000;
   assign mem[329151:329120] = 32'b00000110111111110001010110001000;
   assign mem[329183:329152] = 32'b11011111010000101100100011000000;
   assign mem[329215:329184] = 32'b00000110110100101011110010101000;
   assign mem[329247:329216] = 32'b11111010011111010001010111110000;
   assign mem[329279:329248] = 32'b00000001100000011011001000101010;
   assign mem[329311:329280] = 32'b00000100110111110101111011010000;
   assign mem[329343:329312] = 32'b11111110100000010111110110111000;
   assign mem[329375:329344] = 32'b00000101110110111010011110101000;
   assign mem[329407:329376] = 32'b11110000001101010101001110110000;
   assign mem[329439:329408] = 32'b00000111100100110000100110111000;
   assign mem[329471:329440] = 32'b11111001111000111001110010010000;
   assign mem[329503:329472] = 32'b11111101101110000000011011110100;
   assign mem[329535:329504] = 32'b11111100010001111101110100110000;
   assign mem[329567:329536] = 32'b00000011110010101001011011000000;
   assign mem[329599:329568] = 32'b00000001011100111000011101001000;
   assign mem[329631:329600] = 32'b11111001100101101111111101000000;
   assign mem[329663:329632] = 32'b00001001111110000111000011010000;
   assign mem[329695:329664] = 32'b00000011001001011101110111110100;
   assign mem[329727:329696] = 32'b11111110010001110100101000001110;
   assign mem[329759:329728] = 32'b11110010010010010111000110110000;
   assign mem[329791:329760] = 32'b11111100100001010110001110101100;
   assign mem[329823:329792] = 32'b11111011000000101001000100000000;
   assign mem[329855:329824] = 32'b00001011110111111101010101110000;
   assign mem[329887:329856] = 32'b11111101110000100111101110100000;
   assign mem[329919:329888] = 32'b11110011111110101101010110110000;
   assign mem[329951:329920] = 32'b00000100001110101111001000100000;
   assign mem[329983:329952] = 32'b00000110011000000111100100000000;
   assign mem[330015:329984] = 32'b00000000100011111111011010110110;
   assign mem[330047:330016] = 32'b11111101010011100111110010110100;
   assign mem[330079:330048] = 32'b00000000010100110110110111000001;
   assign mem[330111:330080] = 32'b11111011000100101010001001100000;
   assign mem[330143:330112] = 32'b00000000100100110110010011100011;
   assign mem[330175:330144] = 32'b00001000001001001000110001100000;
   assign mem[330207:330176] = 32'b00001011100001110100101000010000;
   assign mem[330239:330208] = 32'b11100110011110101001010010000000;
   assign mem[330271:330240] = 32'b11101000100110000101001110100000;
   assign mem[330303:330272] = 32'b00000101010110010111001001111000;
   assign mem[330335:330304] = 32'b11111010110101001011011001101000;
   assign mem[330367:330336] = 32'b00001000110100010110101000000000;
   assign mem[330399:330368] = 32'b11111110110000111001001001000000;
   assign mem[330431:330400] = 32'b00000101010010011011000101100000;
   assign mem[330463:330432] = 32'b11100001100001001101011111100000;
   assign mem[330495:330464] = 32'b00000010001000000011100110011100;
   assign mem[330527:330496] = 32'b11110101100111000110111111100000;
   assign mem[330559:330528] = 32'b00000010011100111100010010001000;
   assign mem[330591:330560] = 32'b00000101111100101110100010000000;
   assign mem[330623:330592] = 32'b00000100010001010000111010001000;
   assign mem[330655:330624] = 32'b00000110000000011111000100111000;
   assign mem[330687:330656] = 32'b11110100101111110011000011010000;
   assign mem[330719:330688] = 32'b11111010001010011111010110010000;
   assign mem[330751:330720] = 32'b11111010101110001000100000110000;
   assign mem[330783:330752] = 32'b11111111011010011000100000001011;
   assign mem[330815:330784] = 32'b11111001101001010010110000010000;
   assign mem[330847:330816] = 32'b00000001110000010111011000100110;
   assign mem[330879:330848] = 32'b11111001111100100111000101001000;
   assign mem[330911:330880] = 32'b00000000000000111111011111011101;
   assign mem[330943:330912] = 32'b00001001011010111100001000110000;
   assign mem[330975:330944] = 32'b11111100010011100011111000110000;
   assign mem[331007:330976] = 32'b11111011111011111001000111001000;
   assign mem[331039:331008] = 32'b11111001000000011011001100110000;
   assign mem[331071:331040] = 32'b11111001110011001110011101010000;
   assign mem[331103:331072] = 32'b00000001111001011101011000001100;
   assign mem[331135:331104] = 32'b00000111011100001011000010001000;
   assign mem[331167:331136] = 32'b00000011000100000000001000011000;
   assign mem[331199:331168] = 32'b11111010010100011111111101110000;
   assign mem[331231:331200] = 32'b11111111011010001011011010010001;
   assign mem[331263:331232] = 32'b11110100111000001100011001100000;
   assign mem[331295:331264] = 32'b11110011111100111010011000000000;
   assign mem[331327:331296] = 32'b11111011000011001000000101001000;
   assign mem[331359:331328] = 32'b00000001110110000111011101101000;
   assign mem[331391:331360] = 32'b00000000000110000111000001111000;
   assign mem[331423:331392] = 32'b00000010010101111101001110010000;
   assign mem[331455:331424] = 32'b00000100100011111000110100110000;
   assign mem[331487:331456] = 32'b00000000001010011011000111111101;
   assign mem[331519:331488] = 32'b00001000001000000001100111010000;
   assign mem[331551:331520] = 32'b00000011001100100111101111110000;
   assign mem[331583:331552] = 32'b00000100111100011010011101101000;
   assign mem[331615:331584] = 32'b11111010010110110010010101011000;
   assign mem[331647:331616] = 32'b11110111111110101011010000000000;
   assign mem[331679:331648] = 32'b00000001111010111111000010100000;
   assign mem[331711:331680] = 32'b11111100000001100111100100011000;
   assign mem[331743:331712] = 32'b11111111111111110011111111100100;
   assign mem[331775:331744] = 32'b11111101000110000001101110110000;
   assign mem[331807:331776] = 32'b11111111110000000010011001110110;
   assign mem[331839:331808] = 32'b00001100011110000111011101110000;
   assign mem[331871:331840] = 32'b00000001111010011001000000101000;
   assign mem[331903:331872] = 32'b00001010101101011101100011110000;
   assign mem[331935:331904] = 32'b11111010011100111011001010001000;
   assign mem[331967:331936] = 32'b00000001000100001111000000011010;
   assign mem[331999:331968] = 32'b00000010010111110000111111100000;
   assign mem[332031:332000] = 32'b00000011101110110010010110101100;
   assign mem[332063:332032] = 32'b11111101111101010110001110000000;
   assign mem[332095:332064] = 32'b00000000110001100110010001000110;
   assign mem[332127:332096] = 32'b11111011110100110010010001010000;
   assign mem[332159:332128] = 32'b00000010010010101111000111110100;
   assign mem[332191:332160] = 32'b00000010111110101010011010000000;
   assign mem[332223:332192] = 32'b00000001011001001011000110101100;
   assign mem[332255:332224] = 32'b11111111110000101010101011101010;
   assign mem[332287:332256] = 32'b11111001001110111110001000101000;
   assign mem[332319:332288] = 32'b00000101001100110100010011110000;
   assign mem[332351:332320] = 32'b00000001011101101101001000010010;
   assign mem[332383:332352] = 32'b00000000011011001011110101100001;
   assign mem[332415:332384] = 32'b11110000001100110010101011010000;
   assign mem[332447:332416] = 32'b00000010100110010101110110010100;
   assign mem[332479:332448] = 32'b00000110100101110111000111110000;
   assign mem[332511:332480] = 32'b00000001111101110011001011111010;
   assign mem[332543:332512] = 32'b00000001011110101110111011101110;
   assign mem[332575:332544] = 32'b00000011011101010001011011000000;
   assign mem[332607:332576] = 32'b11111110011101111100011011010010;
   assign mem[332639:332608] = 32'b00000100000110001100010111101000;
   assign mem[332671:332640] = 32'b11111011011010010011110010011000;
   assign mem[332703:332672] = 32'b00000000100010101110100110011111;
   assign mem[332735:332704] = 32'b11111100101011001100100001100000;
   assign mem[332767:332736] = 32'b00000111100011110001011001000000;
   assign mem[332799:332768] = 32'b11111001000000111010111000101000;
   assign mem[332831:332800] = 32'b11111111010001001010101001010111;
   assign mem[332863:332832] = 32'b00000000010111110110010000101101;
   assign mem[332895:332864] = 32'b00000101000101001110000001111000;
   assign mem[332927:332896] = 32'b11111101111011001001100111111000;
   assign mem[332959:332928] = 32'b11111111110010101101101001110001;
   assign mem[332991:332960] = 32'b00000000010010011111110110011101;
   assign mem[333023:332992] = 32'b11111101111010101000101111011100;
   assign mem[333055:333024] = 32'b11111100101011100111011011110000;
   assign mem[333087:333056] = 32'b11110101111111111010110001000000;
   assign mem[333119:333088] = 32'b00000010011100110001000101111100;
   assign mem[333151:333120] = 32'b00000110001101111100100000111000;
   assign mem[333183:333152] = 32'b11111010111101110101011010111000;
   assign mem[333215:333184] = 32'b00000000000110011010100010111011;
   assign mem[333247:333216] = 32'b11110111110101000001010101100000;
   assign mem[333279:333248] = 32'b11111110110101010001101111100000;
   assign mem[333311:333280] = 32'b11110111000101010101100100000000;
   assign mem[333343:333312] = 32'b00000100001100110101011011001000;
   assign mem[333375:333344] = 32'b11111100010010100001011001010100;
   assign mem[333407:333376] = 32'b11111111100100000110010000111100;
   assign mem[333439:333408] = 32'b00000000110001100110110110000010;
   assign mem[333471:333440] = 32'b11111011010100111101000101110000;
   assign mem[333503:333472] = 32'b00000000000000000001001100110110;
   assign mem[333535:333504] = 32'b11111001011100001111100111000000;
   assign mem[333567:333536] = 32'b00000010011000110001001101011100;
   assign mem[333599:333568] = 32'b00001010100011101101000001110000;
   assign mem[333631:333600] = 32'b00000100001000110000101011001000;
   assign mem[333663:333632] = 32'b11110100100110011111000011010000;
   assign mem[333695:333664] = 32'b11111011111000010011101110101000;
   assign mem[333727:333696] = 32'b11111001110001111100110110101000;
   assign mem[333759:333728] = 32'b00000000001000001001001010011101;
   assign mem[333791:333760] = 32'b11111110010101001011001000000010;
   assign mem[333823:333792] = 32'b00000011100011100111111101001000;
   assign mem[333855:333824] = 32'b00000100101110100101111011000000;
   assign mem[333887:333856] = 32'b11111111000110111100110111000000;
   assign mem[333919:333888] = 32'b00000100011111110001001110010000;
   assign mem[333951:333920] = 32'b00000001010001100101010011001000;
   assign mem[333983:333952] = 32'b11110100111000000110101011010000;
   assign mem[334015:333984] = 32'b00000001111110110000111111111010;
   assign mem[334047:334016] = 32'b00000011101001101110011000011100;
   assign mem[334079:334048] = 32'b11111101010111001111101110110100;
   assign mem[334111:334080] = 32'b00000100001000000111001001011000;
   assign mem[334143:334112] = 32'b00000010011010100000100010100000;
   assign mem[334175:334144] = 32'b00000011001100011001010111100100;
   assign mem[334207:334176] = 32'b11110101001001110010010001110000;
   assign mem[334239:334208] = 32'b00000000100100011010001101001100;
   assign mem[334271:334240] = 32'b11111100010001010011010101110100;
   assign mem[334303:334272] = 32'b00000110010011010110010100000000;
   assign mem[334335:334304] = 32'b11111110011001100011011110001000;
   assign mem[334367:334336] = 32'b00000001110000011110010111010100;
   assign mem[334399:334368] = 32'b11111000111100111110111001001000;
   assign mem[334431:334400] = 32'b11111111101101110111011010111110;
   assign mem[334463:334432] = 32'b11111110101101100000100011110000;
   assign mem[334495:334464] = 32'b00000101010011010011111111100000;
   assign mem[334527:334496] = 32'b11111110000001001011011111110010;
   assign mem[334559:334528] = 32'b00000000110110110110010011111100;
   assign mem[334591:334560] = 32'b11111011111011010110110001111000;
   assign mem[334623:334592] = 32'b11111000011111101111010000100000;
   assign mem[334655:334624] = 32'b00000001100010111110011100010100;
   assign mem[334687:334656] = 32'b11111101110011000111000100011000;
   assign mem[334719:334688] = 32'b00000011001011100001010001011100;
   assign mem[334751:334720] = 32'b00000100010011001000001000010000;
   assign mem[334783:334752] = 32'b00000100000001000110100010001000;
   assign mem[334815:334784] = 32'b00000100100110111001110101001000;
   assign mem[334847:334816] = 32'b11110100010010001100101001100000;
   assign mem[334879:334848] = 32'b00000100110011110110111011111000;
   assign mem[334911:334880] = 32'b11111101010111000010001110001100;
   assign mem[334943:334912] = 32'b00000001000001011110110111001000;
   assign mem[334975:334944] = 32'b11110110110100111011001111110000;
   assign mem[335007:334976] = 32'b00001000100011100001110001110000;
   assign mem[335039:335008] = 32'b11111000110010101000011101100000;
   assign mem[335071:335040] = 32'b00000100011110111011001011110000;
   assign mem[335103:335072] = 32'b11110100011100110110011010010000;
   assign mem[335135:335104] = 32'b00000010111110011101011010111100;
   assign mem[335167:335136] = 32'b11111111111100010110010101101101;
   assign mem[335199:335168] = 32'b00000001111101101100010110010110;
   assign mem[335231:335200] = 32'b11111011001110110110110001000000;
   assign mem[335263:335232] = 32'b00000101000100111111101101011000;
   assign mem[335295:335264] = 32'b11111011000101000000011000001000;
   assign mem[335327:335296] = 32'b00000001111100001101111101010000;
   assign mem[335359:335328] = 32'b11111111110100111111000000110101;
   assign mem[335391:335360] = 32'b00000001100011100010011001000110;
   assign mem[335423:335392] = 32'b11110011000011011110001011110000;
   assign mem[335455:335424] = 32'b11111111111010011110001001110101;
   assign mem[335487:335456] = 32'b11111001111100000110001010010000;
   assign mem[335519:335488] = 32'b11111110001111001110000111001100;
   assign mem[335551:335520] = 32'b00000001001100011111101101101000;
   assign mem[335583:335552] = 32'b11111110001101110010101001000100;
   assign mem[335615:335584] = 32'b11111001100100110110100111111000;
   assign mem[335647:335616] = 32'b00000110000001111011111001111000;
   assign mem[335679:335648] = 32'b00000100001101101110110100111000;
   assign mem[335711:335680] = 32'b00000100011011110001101101101000;
   assign mem[335743:335712] = 32'b11111101000111111001010001000000;
   assign mem[335775:335744] = 32'b11110111100111000111100110100000;
   assign mem[335807:335776] = 32'b11110101101001011000011010000000;
   assign mem[335839:335808] = 32'b00000111001111100111101011101000;
   assign mem[335871:335840] = 32'b11111000110111111100000000100000;
   assign mem[335903:335872] = 32'b11111011001111000101001011100000;
   assign mem[335935:335904] = 32'b00010011000001110001101001000000;
   assign mem[335967:335936] = 32'b11111111011111010010011100010001;
   assign mem[335999:335968] = 32'b11110111010011110110110100000000;
   assign mem[336031:336000] = 32'b00000010110101011000000101111000;
   assign mem[336063:336032] = 32'b00000100000001101011110001110000;
   assign mem[336095:336064] = 32'b11111001010100000011110111111000;
   assign mem[336127:336096] = 32'b11110111111110011110100010110000;
   assign mem[336159:336128] = 32'b11111110110011011101100111111000;
   assign mem[336191:336160] = 32'b11110101001100100001110101000000;
   assign mem[336223:336192] = 32'b00000101010110111101011000000000;
   assign mem[336255:336224] = 32'b00000100000000010011110001010000;
   assign mem[336287:336256] = 32'b00000001000101101000110010110100;
   assign mem[336319:336288] = 32'b00000111111011101010011001000000;
   assign mem[336351:336320] = 32'b11111001001011001011001110010000;
   assign mem[336383:336352] = 32'b00000011100110101100101000110000;
   assign mem[336415:336384] = 32'b00000111000010000110110000011000;
   assign mem[336447:336416] = 32'b11111111001000000100011000010000;
   assign mem[336479:336448] = 32'b11111001010111001000000011011000;
   assign mem[336511:336480] = 32'b11110110011100110001000111110000;
   assign mem[336543:336512] = 32'b11110100111010001101110100110000;
   assign mem[336575:336544] = 32'b00000110100101101110010100000000;
   assign mem[336607:336576] = 32'b00001000000100111101011001000000;
   assign mem[336639:336608] = 32'b00000000111111011100001111101111;
   assign mem[336671:336640] = 32'b00000010100001101010111101000100;
   assign mem[336703:336672] = 32'b00000010110111011001101011100000;
   assign mem[336735:336704] = 32'b00000011011011001110100111100100;
   assign mem[336767:336736] = 32'b11111000100000101110111010110000;
   assign mem[336799:336768] = 32'b00000010010101000101101101110000;
   assign mem[336831:336800] = 32'b11111100100010101010001011000100;
   assign mem[336863:336832] = 32'b11110111011110100011000101010000;
   assign mem[336895:336864] = 32'b11110101000100101100111110100000;
   assign mem[336927:336896] = 32'b00000001000010000110111111010100;
   assign mem[336959:336928] = 32'b00001000000011111110010010000000;
   assign mem[336991:336960] = 32'b11110010011101111000101011110000;
   assign mem[337023:336992] = 32'b00001000001011010000001011110000;
   assign mem[337055:337024] = 32'b00000001001001000111011010100110;
   assign mem[337087:337056] = 32'b00000011010100111100100001100000;
   assign mem[337119:337088] = 32'b11110011111101011110010011110000;
   assign mem[337151:337120] = 32'b00001000101001110000101100110000;
   assign mem[337183:337152] = 32'b11111001101001001011001011010000;
   assign mem[337215:337184] = 32'b00000110110011000100101010010000;
   assign mem[337247:337216] = 32'b11110011010100110001000000010000;
   assign mem[337279:337248] = 32'b00000000111100101010010101011100;
   assign mem[337311:337280] = 32'b00000000010000110101000000110000;
   assign mem[337343:337312] = 32'b00000000101001000001001110110111;
   assign mem[337375:337344] = 32'b11111101010010000111110110111000;
   assign mem[337407:337376] = 32'b00000001011101010100100100001100;
   assign mem[337439:337408] = 32'b00000101100110100101000011001000;
   assign mem[337471:337440] = 32'b11111011110001000100001011010000;
   assign mem[337503:337472] = 32'b00000010101101001010011110011000;
   assign mem[337535:337504] = 32'b00000000011000000100100111110111;
   assign mem[337567:337536] = 32'b11111010110011110011000101100000;
   assign mem[337599:337568] = 32'b11111110111010100011111000001110;
   assign mem[337631:337600] = 32'b00000001000100000000110101101010;
   assign mem[337663:337632] = 32'b11110111100101001000111100100000;
   assign mem[337695:337664] = 32'b11111011010001101111011010111000;
   assign mem[337727:337696] = 32'b11111100011100010110110011111000;
   assign mem[337759:337728] = 32'b00000100001010100110110011010000;
   assign mem[337791:337760] = 32'b00000010110110011001110100001000;
   assign mem[337823:337792] = 32'b11111001101101110000111001000000;
   assign mem[337855:337824] = 32'b00000001011001001111010000000010;
   assign mem[337887:337856] = 32'b11111011101011100011011111001000;
   assign mem[337919:337888] = 32'b00000011101010011111110110101100;
   assign mem[337951:337920] = 32'b00000110011001100010000100111000;
   assign mem[337983:337952] = 32'b00000101001000110101101101111000;
   assign mem[338015:337984] = 32'b00001000110010101000011010100000;
   assign mem[338047:338016] = 32'b11110011111110000100001110010000;
   assign mem[338079:338048] = 32'b11111101111010110001111011001000;
   assign mem[338111:338080] = 32'b11110101000000111000000011110000;
   assign mem[338143:338112] = 32'b11111111000010000000010110000100;
   assign mem[338175:338144] = 32'b00000000011010100110011000100110;
   assign mem[338207:338176] = 32'b00001011100001011110101001000000;
   assign mem[338239:338208] = 32'b11100111101011010011110001100000;
   assign mem[338271:338240] = 32'b00000100100110110100110001001000;
   assign mem[338303:338272] = 32'b11111101100110000101000001101000;
   assign mem[338335:338304] = 32'b00000100110100000010110011010000;
   assign mem[338367:338336] = 32'b11110100001101100001111010000000;
   assign mem[338399:338368] = 32'b00000110101100001010111001010000;
   assign mem[338431:338400] = 32'b11110110100001110111110100110000;
   assign mem[338463:338432] = 32'b00000111001011100010010100001000;
   assign mem[338495:338464] = 32'b11111100010100101000101111110100;
   assign mem[338527:338496] = 32'b00000100111110111100100111110000;
   assign mem[338559:338528] = 32'b00000001101110111000001101100110;
   assign mem[338591:338560] = 32'b00000010110101001010110100010000;
   assign mem[338623:338592] = 32'b11111101101111010110101010000100;
   assign mem[338655:338624] = 32'b11111101111011100001001111010100;
   assign mem[338687:338656] = 32'b11110110011000011111110011000000;
   assign mem[338719:338688] = 32'b00000100010000110011011000010000;
   assign mem[338751:338720] = 32'b11111100000010111000110101001000;
   assign mem[338783:338752] = 32'b11111000110110110000101111101000;
   assign mem[338815:338784] = 32'b11111110001000111010101111000110;
   assign mem[338847:338816] = 32'b11111110110110000000001000111000;
   assign mem[338879:338848] = 32'b00001000011001001101101000010000;
   assign mem[338911:338880] = 32'b11111001101110011000001100101000;
   assign mem[338943:338912] = 32'b11111111101001010101101000100111;
   assign mem[338975:338944] = 32'b00000101110000011111101110110000;
   assign mem[339007:338976] = 32'b11111011011100010001011110100000;
   assign mem[339039:339008] = 32'b11111000000010100111001111001000;
   assign mem[339071:339040] = 32'b11111001000011111101000100110000;
   assign mem[339103:339072] = 32'b11111100010001100101011010010100;
   assign mem[339135:339104] = 32'b00001011101110111111010000000000;
   assign mem[339167:339136] = 32'b00000010100110001111100010111000;
   assign mem[339199:339168] = 32'b11111000011011100000110000110000;
   assign mem[339231:339200] = 32'b11111101001011100111111000111000;
   assign mem[339263:339232] = 32'b00000011000000001001010011110100;
   assign mem[339295:339264] = 32'b11111000100100101110011101110000;
   assign mem[339327:339296] = 32'b00000101101010110101000111111000;
   assign mem[339359:339328] = 32'b00000110011111100011100000111000;
   assign mem[339391:339360] = 32'b00000101010001000000110000110000;
   assign mem[339423:339392] = 32'b11110101001001010010000100100000;
   assign mem[339455:339424] = 32'b00000000010101010111101110000100;
   assign mem[339487:339456] = 32'b11110111010000011011111101000000;
   assign mem[339519:339488] = 32'b11111111101100101011100110111101;
   assign mem[339551:339520] = 32'b11111101010010101000100011011100;
   assign mem[339583:339552] = 32'b11111110110011001101010000010000;
   assign mem[339615:339584] = 32'b11111100010101101000100100010100;
   assign mem[339647:339616] = 32'b00001000001000100001010111110000;
   assign mem[339679:339648] = 32'b11111111000110000110001011111010;
   assign mem[339711:339680] = 32'b00000101010101010101000101101000;
   assign mem[339743:339712] = 32'b11111110001100101111110111001110;
   assign mem[339775:339744] = 32'b00000101111000011101101011011000;
   assign mem[339807:339776] = 32'b11101110110100010000100110100000;
   assign mem[339839:339808] = 32'b00000011010111100110000000110100;
   assign mem[339871:339840] = 32'b11111101111010111110001010010100;
   assign mem[339903:339872] = 32'b11111100011111110111010110101100;
   assign mem[339935:339904] = 32'b00000001010000001101011111111110;
   assign mem[339967:339936] = 32'b11111001100101001011011111111000;
   assign mem[339999:339968] = 32'b00000011000010011110100100001000;
   assign mem[340031:340000] = 32'b00000010110000111101111111111100;
   assign mem[340063:340032] = 32'b00000010010111000000011000011000;
   assign mem[340095:340064] = 32'b11110010110111001000111101100000;
   assign mem[340127:340096] = 32'b00000000001100000001000000111000;
   assign mem[340159:340128] = 32'b00000111100010011001010111001000;
   assign mem[340191:340160] = 32'b11100100011001101000100001000000;
   assign mem[340223:340192] = 32'b00001000000001111001110000010000;
   assign mem[340255:340224] = 32'b11111110111100011101110011011010;
   assign mem[340287:340256] = 32'b00000000111001100000110010001111;
   assign mem[340319:340288] = 32'b00000011010010011101001010101100;
   assign mem[340351:340320] = 32'b00000110011111111010101111001000;
   assign mem[340383:340352] = 32'b11011111111100000100101100000000;
   assign mem[340415:340384] = 32'b00000011110110111100110010000100;
   assign mem[340447:340416] = 32'b11111000101111010001011011010000;
   assign mem[340479:340448] = 32'b00000001111000000000010100010100;
   assign mem[340511:340480] = 32'b00000101010011011000110110100000;
   assign mem[340543:340512] = 32'b11101110111001010010011011100000;
   assign mem[340575:340544] = 32'b00000001000010010010000100011110;
   assign mem[340607:340576] = 32'b11101111100100100011001110100000;
   assign mem[340639:340608] = 32'b00000011011101001001101100110000;
   assign mem[340671:340640] = 32'b11111100011110010010111011011000;
   assign mem[340703:340672] = 32'b00000101001011000001010010101000;
   assign mem[340735:340704] = 32'b11111100010010100110011101000100;
   assign mem[340767:340736] = 32'b00000001000101001111111110101010;
   assign mem[340799:340768] = 32'b00000110001110110110111010111000;
   assign mem[340831:340800] = 32'b11111011110010110010010000010000;
   assign mem[340863:340832] = 32'b00000000110011110110001110110110;
   assign mem[340895:340864] = 32'b00000101110100111111100001010000;
   assign mem[340927:340896] = 32'b00000010000100010011000010010100;
   assign mem[340959:340928] = 32'b00000010101010111011000000111100;
   assign mem[340991:340960] = 32'b00000101010000011001000100000000;
   assign mem[341023:340992] = 32'b11110111110000111110000000010000;
   assign mem[341055:341024] = 32'b00000011000100010110100001011100;
   assign mem[341087:341056] = 32'b11111100100001001010001001010100;
   assign mem[341119:341088] = 32'b00000011001100001010111111000100;
   assign mem[341151:341120] = 32'b11111001110000101000101100011000;
   assign mem[341183:341152] = 32'b00000001010010110100101101110010;
   assign mem[341215:341184] = 32'b11111001100110110011001100101000;
   assign mem[341247:341216] = 32'b00000110111011110101111011111000;
   assign mem[341279:341248] = 32'b00000100000010011011010100001000;
   assign mem[341311:341280] = 32'b00000011100001110111000101011000;
   assign mem[341343:341312] = 32'b11110100001001111100000010110000;
   assign mem[341375:341344] = 32'b00000100000111101100000110010000;
   assign mem[341407:341376] = 32'b11110111001101100111101110100000;
   assign mem[341439:341408] = 32'b00000101011111100100001101110000;
   assign mem[341471:341440] = 32'b00000000011011101111101100001010;
   assign mem[341503:341472] = 32'b11110100101111100011100001000000;
   assign mem[341535:341504] = 32'b11110100010010101010000010010000;
   assign mem[341567:341536] = 32'b00001101101010110111110101010000;
   assign mem[341599:341568] = 32'b00000000111110000001000010011001;
   assign mem[341631:341600] = 32'b00001000001010010101110000000000;
   assign mem[341663:341632] = 32'b00000010111011100100100010100000;
   assign mem[341695:341664] = 32'b00000001010010010101010011010110;
   assign mem[341727:341696] = 32'b11110100000010101110000000010000;
   assign mem[341759:341728] = 32'b00000001110010011001101110100110;
   assign mem[341791:341760] = 32'b00000001110011111000000100110010;
   assign mem[341823:341792] = 32'b11110100111000100111101110100000;
   assign mem[341855:341824] = 32'b00000011001101100000111010001000;
   assign mem[341887:341856] = 32'b11111011100010111001110100001000;
   assign mem[341919:341888] = 32'b00000100111110011100010111010000;
   assign mem[341951:341920] = 32'b11111110100100000101100110011010;
   assign mem[341983:341952] = 32'b11111110111110110000000110010010;
   assign mem[342015:341984] = 32'b11110011101111110111000110110000;
   assign mem[342047:342016] = 32'b00000011111110000100111101111100;
   assign mem[342079:342048] = 32'b00000001011011001000111111110000;
   assign mem[342111:342080] = 32'b00000000101110010000111110011110;
   assign mem[342143:342112] = 32'b11111000011111111001010000001000;
   assign mem[342175:342144] = 32'b11110011100001110011000000100000;
   assign mem[342207:342176] = 32'b00001000111001100001010101100000;
   assign mem[342239:342208] = 32'b11110110100001011011011111100000;
   assign mem[342271:342240] = 32'b11111001001101100100011011011000;
   assign mem[342303:342272] = 32'b00000100111100000100001111101000;
   assign mem[342335:342304] = 32'b11111101001100110111111000100000;
   assign mem[342367:342336] = 32'b00000100011001000000100000010000;
   assign mem[342399:342368] = 32'b00000001001011000110011100111000;
   assign mem[342431:342400] = 32'b00000101110101111101011110101000;
   assign mem[342463:342432] = 32'b00000011110001010101001011101100;
   assign mem[342495:342464] = 32'b11110101100101011001010011010000;
   assign mem[342527:342496] = 32'b11111000011111101010010111111000;
   assign mem[342559:342528] = 32'b00000100110100111010001111110000;
   assign mem[342591:342560] = 32'b11111000101101011001110111010000;
   assign mem[342623:342592] = 32'b00000011011010101101000101010100;
   assign mem[342655:342624] = 32'b11111010001111011000010101110000;
   assign mem[342687:342656] = 32'b00001001110010000100010010100000;
   assign mem[342719:342688] = 32'b11111111011101010110000101110001;
   assign mem[342751:342720] = 32'b00000010011010100111110000001100;
   assign mem[342783:342752] = 32'b00000001100101100101010010010010;
   assign mem[342815:342784] = 32'b11111110000001001111011010010100;
   assign mem[342847:342816] = 32'b00000011010111100000101111100100;
   assign mem[342879:342848] = 32'b11111101111100110110100011101000;
   assign mem[342911:342880] = 32'b00000011001110101001011010010000;
   assign mem[342943:342912] = 32'b00000011001010101110010110010000;
   assign mem[342975:342944] = 32'b00000010011010100010100001101100;
   assign mem[343007:342976] = 32'b00000011000101001101011010001100;
   assign mem[343039:343008] = 32'b00000000011001001110001110011100;
   assign mem[343071:343040] = 32'b00000001000001110000010000110100;
   assign mem[343103:343072] = 32'b11111001010101111000010000111000;
   assign mem[343135:343104] = 32'b00000110010101111001110011011000;
   assign mem[343167:343136] = 32'b11111101110110110000101101000100;
   assign mem[343199:343168] = 32'b00000100000010011101110001011000;
   assign mem[343231:343200] = 32'b11111001000110001011001101110000;
   assign mem[343263:343232] = 32'b00000011001110001110000100100000;
   assign mem[343295:343264] = 32'b11111100001010111001101101010100;
   assign mem[343327:343296] = 32'b00000101110110100011101001101000;
   assign mem[343359:343328] = 32'b11111111111011100000100110000001;
   assign mem[343391:343360] = 32'b11111111000111101001010111001100;
   assign mem[343423:343392] = 32'b00000100010001001001111110011000;
   assign mem[343455:343424] = 32'b00000110000001000011101111110000;
   assign mem[343487:343456] = 32'b11110100010100100100100000010000;
   assign mem[343519:343488] = 32'b11110111110111011100101010000000;
   assign mem[343551:343520] = 32'b11110011110100000001000111110000;
   assign mem[343583:343552] = 32'b11111111011110001000000001101100;
   assign mem[343615:343584] = 32'b00000000011010001000101110010110;
   assign mem[343647:343616] = 32'b00001000010101100010111000010000;
   assign mem[343679:343648] = 32'b11111011100111000100010010011000;
   assign mem[343711:343680] = 32'b00000000001001001100000001011010;
   assign mem[343743:343712] = 32'b11111000001110001111101000010000;
   assign mem[343775:343744] = 32'b00000101110010011100010011001000;
   assign mem[343807:343776] = 32'b11110000001101110010101001000000;
   assign mem[343839:343808] = 32'b00000011001111101001011100011100;
   assign mem[343871:343840] = 32'b11111011111001011101110111000000;
   assign mem[343903:343872] = 32'b11111000000010111100000111010000;
   assign mem[343935:343904] = 32'b00000010101011111110101000010100;
   assign mem[343967:343936] = 32'b00001001100110110001100111110000;
   assign mem[343999:343968] = 32'b11111010000001010000001011000000;
   assign mem[344031:344000] = 32'b00000011011110101011000001100100;
   assign mem[344063:344032] = 32'b00000001011111000011110100000010;
   assign mem[344095:344064] = 32'b11111100110000101000101000100000;
   assign mem[344127:344096] = 32'b00001111011110110010100000100000;
   assign mem[344159:344128] = 32'b11111010000011100001011101011000;
   assign mem[344191:344160] = 32'b00000100001111110001010101110000;
   assign mem[344223:344192] = 32'b11111110010001000111101001101010;
   assign mem[344255:344224] = 32'b11111010110111000010011110101000;
   assign mem[344287:344256] = 32'b00000000010000001011101001011111;
   assign mem[344319:344288] = 32'b11111111101010011011100000010111;
   assign mem[344351:344320] = 32'b11111110010110010001011000011010;
   assign mem[344383:344352] = 32'b11111111011101110000010010011000;
   assign mem[344415:344384] = 32'b00000000011010001010000011010000;
   assign mem[344447:344416] = 32'b11111111110010001111000001110111;
   assign mem[344479:344448] = 32'b00000001011101111110100001000010;
   assign mem[344511:344480] = 32'b11111111100100100010110101011011;
   assign mem[344543:344512] = 32'b11111101110010001001000101111000;
   assign mem[344575:344544] = 32'b11111100011001000100111110101000;
   assign mem[344607:344576] = 32'b11111011101100000101000001101000;
   assign mem[344639:344608] = 32'b00000011001111010100100101011100;
   assign mem[344671:344640] = 32'b00000000100111001011101111111110;
   assign mem[344703:344672] = 32'b00000010100101110001010100010100;
   assign mem[344735:344704] = 32'b11111110101010111111110011001110;
   assign mem[344767:344736] = 32'b11111100110111111110101001001000;
   assign mem[344799:344768] = 32'b00001011000010011000100010000000;
   assign mem[344831:344800] = 32'b11111110011100100111100100001100;
   assign mem[344863:344832] = 32'b11111001110010110010001010010000;
   assign mem[344895:344864] = 32'b00000010111110010111000011010000;
   assign mem[344927:344896] = 32'b11111011001000010010010001100000;
   assign mem[344959:344928] = 32'b00000100001110100110110111100000;
   assign mem[344991:344960] = 32'b11111111111010111110011100111111;
   assign mem[345023:344992] = 32'b11111110011100100101110110011000;
   assign mem[345055:345024] = 32'b00000001001000001010111100011010;
   assign mem[345087:345056] = 32'b11111010110001011100100011001000;
   assign mem[345119:345088] = 32'b00000100001010001000100100010000;
   assign mem[345151:345120] = 32'b00000011000110000110010101010100;
   assign mem[345183:345152] = 32'b11111110101111110010001010101110;
   assign mem[345215:345184] = 32'b00000001110110111010100110111000;
   assign mem[345247:345216] = 32'b11111100010001110110011011110100;
   assign mem[345279:345248] = 32'b00000000111110101000100111111110;
   assign mem[345311:345280] = 32'b00000111001101111110001100000000;
   assign mem[345343:345312] = 32'b00000011110111000001010001110100;
   assign mem[345375:345344] = 32'b11111010110100101110111001111000;
   assign mem[345407:345376] = 32'b11110111000110010110110110100000;
   assign mem[345439:345408] = 32'b11111011000111000010010111010000;
   assign mem[345471:345440] = 32'b11111010011010101011010001111000;
   assign mem[345503:345472] = 32'b00000110011000010011100101111000;
   assign mem[345535:345504] = 32'b11111110100001111101101010101100;
   assign mem[345567:345536] = 32'b00000000011010111101011110011101;
   assign mem[345599:345568] = 32'b11111011001101000101111010001000;
   assign mem[345631:345600] = 32'b11111110111100000001001100010100;
   assign mem[345663:345632] = 32'b11111010101010110100101101110000;
   assign mem[345695:345664] = 32'b00000110000101101001000111100000;
   assign mem[345727:345696] = 32'b00000010001011110001100011100100;
   assign mem[345759:345728] = 32'b11111111101110011011011101101100;
   assign mem[345791:345760] = 32'b11111110010101101111011000010110;
   assign mem[345823:345792] = 32'b11111101011101001011101000010100;
   assign mem[345855:345824] = 32'b00000100110110110111010101111000;
   assign mem[345887:345856] = 32'b00000011101011001110111010111000;
   assign mem[345919:345888] = 32'b11111001101011100111100100111000;
   assign mem[345951:345920] = 32'b11111010110011101111011010010000;
   assign mem[345983:345952] = 32'b11110000111000010011100101010000;
   assign mem[346015:345984] = 32'b11110000010000000110010101110000;
   assign mem[346047:346016] = 32'b11111101011000011010011011110000;
   assign mem[346079:346048] = 32'b00000100101011000001101010011000;
   assign mem[346111:346080] = 32'b00000001000110000101011101000010;
   assign mem[346143:346112] = 32'b11111111101111011110101011110101;
   assign mem[346175:346144] = 32'b11111101001011000111101110011000;
   assign mem[346207:346176] = 32'b00000011110110100001100010111100;
   assign mem[346239:346208] = 32'b00000110001010110001111011110000;
   assign mem[346271:346240] = 32'b11111111011111111100100110010100;
   assign mem[346303:346272] = 32'b00000101000001001000111000011000;
   assign mem[346335:346304] = 32'b00000000111001000101011000101000;
   assign mem[346367:346336] = 32'b00001000010010011001001011010000;
   assign mem[346399:346368] = 32'b11111010010000011101011010001000;
   assign mem[346431:346400] = 32'b00001001111100011001100011110000;
   assign mem[346463:346432] = 32'b11110110010000100101011000110000;
   assign mem[346495:346464] = 32'b00000010010011010001001000010100;
   assign mem[346527:346496] = 32'b11101110001001111101010101000000;
   assign mem[346559:346528] = 32'b11111110110111001111001101010110;
   assign mem[346591:346560] = 32'b11111101101101000111111010000100;
   assign mem[346623:346592] = 32'b00000001001001001000000000101100;
   assign mem[346655:346624] = 32'b00000001010000100100111000101000;
   assign mem[346687:346656] = 32'b00001010010100000110000110100000;
   assign mem[346719:346688] = 32'b11110111110101011001100011110000;
   assign mem[346751:346720] = 32'b00000011101101111011011000000100;
   assign mem[346783:346752] = 32'b11111111101011011101110110110000;
   assign mem[346815:346784] = 32'b11111100101110111111011001110000;
   assign mem[346847:346816] = 32'b00000001000011110011101100011010;
   assign mem[346879:346848] = 32'b11111100110011100000111110100100;
   assign mem[346911:346880] = 32'b11110011101010101101001010000000;
   assign mem[346943:346912] = 32'b11111111110110001101010111110110;
   assign mem[346975:346944] = 32'b00000011101010010000001000100000;
   assign mem[347007:346976] = 32'b11111111001001101111000100001100;
   assign mem[347039:347008] = 32'b11111100011011111110111111110000;
   assign mem[347071:347040] = 32'b00000010001110000100101101100000;
   assign mem[347103:347072] = 32'b11101111001010100101110110100000;
   assign mem[347135:347104] = 32'b00000101101001101001010010001000;
   assign mem[347167:347136] = 32'b11111101010110110000000011000100;
   assign mem[347199:347168] = 32'b00000000000110100011011100111010;
   assign mem[347231:347200] = 32'b00000110001001000010110111011000;
   assign mem[347263:347232] = 32'b00000011001011010000111101010100;
   assign mem[347295:347264] = 32'b00001000001001001110000010110000;
   assign mem[347327:347296] = 32'b11111010100011010000101101101000;
   assign mem[347359:347328] = 32'b11111001011100011001001101000000;
   assign mem[347391:347360] = 32'b11110100000010011000100000010000;
   assign mem[347423:347392] = 32'b00000001010111010001100001100000;
   assign mem[347455:347424] = 32'b00000000110001101011001110101001;
   assign mem[347487:347456] = 32'b00001000011100101001101001100000;
   assign mem[347519:347488] = 32'b11111101011101110001110100010100;
   assign mem[347551:347520] = 32'b00000100000010011000111110000000;
   assign mem[347583:347552] = 32'b11111111001010110101101110011110;
   assign mem[347615:347584] = 32'b00000101111111110100101011101000;
   assign mem[347647:347616] = 32'b11111101101100100011110101000100;
   assign mem[347679:347648] = 32'b00000000001010111011101001010001;
   assign mem[347711:347680] = 32'b11111101000100011011000001101100;
   assign mem[347743:347712] = 32'b00000011011001000111110100011000;
   assign mem[347775:347744] = 32'b11110110000100010011010010110000;
   assign mem[347807:347776] = 32'b11111111011100101011101001111110;
   assign mem[347839:347808] = 32'b00000010110010011011110000000000;
   assign mem[347871:347840] = 32'b00000100000000111101011100100000;
   assign mem[347903:347872] = 32'b00000010111101110010011100011100;
   assign mem[347935:347904] = 32'b00000111100100100010101110010000;
   assign mem[347967:347936] = 32'b11110100101010000011101100010000;
   assign mem[347999:347968] = 32'b00000001001010010010101011100110;
   assign mem[348031:348000] = 32'b11111100000001000100000011010000;
   assign mem[348063:348032] = 32'b00000010101101011000011000111100;
   assign mem[348095:348064] = 32'b11111010101111011000000001000000;
   assign mem[348127:348096] = 32'b00001000000110111110110100000000;
   assign mem[348159:348128] = 32'b11111011001011111000011000000000;
   assign mem[348191:348160] = 32'b11111010110001000100000001101000;
   assign mem[348223:348192] = 32'b00000000100001010010010001011001;
   assign mem[348255:348224] = 32'b00000100010001001101101010001000;
   assign mem[348287:348256] = 32'b00000111011001100111110011011000;
   assign mem[348319:348288] = 32'b11111111000010011101000011111100;
   assign mem[348351:348320] = 32'b00000011000010101001000110101100;
   assign mem[348383:348352] = 32'b11111111010110111001100000101011;
   assign mem[348415:348384] = 32'b11110010100110010111010101100000;
   assign mem[348447:348416] = 32'b00000100001111101001101110010000;
   assign mem[348479:348448] = 32'b11111111011000101100101010001110;
   assign mem[348511:348480] = 32'b00010001000111011100111110100000;
   assign mem[348543:348512] = 32'b00000101001110100111000101110000;
   assign mem[348575:348544] = 32'b11101011110011011010110111000000;
   assign mem[348607:348576] = 32'b00001000010010000100010010100000;
   assign mem[348639:348608] = 32'b11111010100010101011111001010000;
   assign mem[348671:348640] = 32'b00001010110001100100010001010000;
   assign mem[348703:348672] = 32'b11111001010101110010000001000000;
   assign mem[348735:348704] = 32'b00001111100110101011001110100000;
   assign mem[348767:348736] = 32'b11100011111111010010001101100000;
   assign mem[348799:348768] = 32'b11111000110110101000001011000000;
   assign mem[348831:348800] = 32'b11111110100010010100110101000010;
   assign mem[348863:348832] = 32'b11110000001100010100100010100000;
   assign mem[348895:348864] = 32'b00000100001101111000001111100000;
   assign mem[348927:348896] = 32'b00000000111111100101011001001111;
   assign mem[348959:348928] = 32'b00000011001001101111010010010100;
   assign mem[348991:348960] = 32'b00000001010011100110010011111010;
   assign mem[349023:348992] = 32'b00000001110000110100010010011000;
   assign mem[349055:349024] = 32'b11101101000111100001010101000000;
   assign mem[349087:349056] = 32'b00000010101101110010111011011000;
   assign mem[349119:349088] = 32'b00000000111101110011110010011010;
   assign mem[349151:349120] = 32'b11110011001011100011000110010000;
   assign mem[349183:349152] = 32'b11100110101010101100010110000000;
   assign mem[349215:349184] = 32'b00000001010110111110010011001100;
   assign mem[349247:349216] = 32'b00000000010001001001110100011000;
   assign mem[349279:349248] = 32'b00000111100111111101000010100000;
   assign mem[349311:349280] = 32'b00000000100110010110010101001110;
   assign mem[349343:349312] = 32'b11110011001000100101100000010000;
   assign mem[349375:349344] = 32'b11111011010010101111100000101000;
   assign mem[349407:349376] = 32'b11111011010110010011011000011000;
   assign mem[349439:349408] = 32'b00001010111010111011010101000000;
   assign mem[349471:349440] = 32'b11110101011001001011010000100000;
   assign mem[349503:349472] = 32'b11111101101010000110001110101100;
   assign mem[349535:349504] = 32'b11111100110010110111110101110100;
   assign mem[349567:349536] = 32'b00000010000011101001111010101100;
   assign mem[349599:349568] = 32'b00000101111010001010111110001000;
   assign mem[349631:349600] = 32'b00000000010100100000010111101011;
   assign mem[349663:349632] = 32'b11110011110010001001110110010000;
   assign mem[349695:349664] = 32'b11111010011111001110000000010000;
   assign mem[349727:349696] = 32'b11111001001011000110100111101000;
   assign mem[349759:349728] = 32'b00000111000101101110101111111000;
   assign mem[349791:349760] = 32'b00000001010010001110001000111010;
   assign mem[349823:349792] = 32'b00000010011111001001111000010100;
   assign mem[349855:349824] = 32'b00000000000001000011101100001011;
   assign mem[349887:349856] = 32'b11111010101111110111100011110000;
   assign mem[349919:349888] = 32'b00000111001100011011001101100000;
   assign mem[349951:349920] = 32'b11110111011001110101101000010000;
   assign mem[349983:349952] = 32'b00000100111010011100011100011000;
   assign mem[350015:349984] = 32'b11111100101000011011001011111100;
   assign mem[350047:350016] = 32'b00000100100110110101110010111000;
   assign mem[350079:350048] = 32'b11111101010010010001111001111100;
   assign mem[350111:350080] = 32'b00000101100011111011011011110000;
   assign mem[350143:350112] = 32'b00010000111100100100010100000000;
   assign mem[350175:350144] = 32'b11111100101111100101010111111000;
   assign mem[350207:350176] = 32'b11110110111011001010100011010000;
   assign mem[350239:350208] = 32'b11110111111000111001110100000000;
   assign mem[350271:350240] = 32'b00000001111010001011110111100100;
   assign mem[350303:350272] = 32'b11110110111101101101110111010000;
   assign mem[350335:350304] = 32'b00001100110010001000111011010000;
   assign mem[350367:350336] = 32'b11111100100001011011011110111100;
   assign mem[350399:350368] = 32'b11110111001010111001111110010000;
   assign mem[350431:350400] = 32'b00000000011101010011000011010011;
   assign mem[350463:350432] = 32'b00000000101110101101101011000010;
   assign mem[350495:350464] = 32'b00000011100011110011000010000100;
   assign mem[350527:350496] = 32'b11111110011101001011101100101000;
   assign mem[350559:350528] = 32'b11111011010010011010010010010000;
   assign mem[350591:350560] = 32'b11111100011011000100100100110100;
   assign mem[350623:350592] = 32'b11111000011111101011001010101000;
   assign mem[350655:350624] = 32'b11111111001101011100101001010110;
   assign mem[350687:350656] = 32'b11111111000001010010011111011111;
   assign mem[350719:350688] = 32'b00001000110001101110111110010000;
   assign mem[350751:350720] = 32'b00000001001110111011101011101110;
   assign mem[350783:350752] = 32'b00001011100000001100010010000000;
   assign mem[350815:350784] = 32'b11111000011011101101110000010000;
   assign mem[350847:350816] = 32'b00001000010011111011001111010000;
   assign mem[350879:350848] = 32'b11111011100011010001111100101000;
   assign mem[350911:350880] = 32'b11111110111111110100111101110000;
   assign mem[350943:350912] = 32'b11110101011111100010010100000000;
   assign mem[350975:350944] = 32'b00000100010011100001110101110000;
   assign mem[351007:350976] = 32'b11101001010000110110011110100000;
   assign mem[351039:351008] = 32'b11111110101000110110101001000110;
   assign mem[351071:351040] = 32'b00000100011011100000110001101000;
   assign mem[351103:351072] = 32'b00000100011100000010110100110000;
   assign mem[351135:351104] = 32'b11111100110010011100001100110000;
   assign mem[351167:351136] = 32'b11111010110111000001101010101000;
   assign mem[351199:351168] = 32'b11111111011100110001101100001001;
   assign mem[351231:351200] = 32'b00000010110000100011000101101000;
   assign mem[351263:351232] = 32'b11111000110000001111010011111000;
   assign mem[351295:351264] = 32'b00000011111001000111111100010000;
   assign mem[351327:351296] = 32'b11111011100110101111011101011000;
   assign mem[351359:351328] = 32'b00000000110011111010100001001011;
   assign mem[351391:351360] = 32'b11111100110110110110001010011000;
   assign mem[351423:351392] = 32'b00000000101011100001111001110010;
   assign mem[351455:351424] = 32'b11111101100101000000010101111000;
   assign mem[351487:351456] = 32'b11111101011011000111100000000000;
   assign mem[351519:351488] = 32'b00000100101110000011110110101000;
   assign mem[351551:351520] = 32'b00000000000100010011001100010010;
   assign mem[351583:351552] = 32'b11111010000111011100001010100000;
   assign mem[351615:351584] = 32'b11111101010111100110010100100100;
   assign mem[351647:351616] = 32'b00000001100011000011110000110010;
   assign mem[351679:351648] = 32'b00000111001110100110111100011000;
   assign mem[351711:351680] = 32'b00000010101100101100111101000100;
   assign mem[351743:351712] = 32'b00000101111001001100001110000000;
   assign mem[351775:351744] = 32'b00000000010011111000001101011000;
   assign mem[351807:351776] = 32'b00000111101001100001100000011000;
   assign mem[351839:351808] = 32'b11111101111000101010011001011000;
   assign mem[351871:351840] = 32'b00000001001011101010010100011100;
   assign mem[351903:351872] = 32'b11111101011011010111111101001000;
   assign mem[351935:351904] = 32'b11111101001001000111111110000000;
   assign mem[351967:351936] = 32'b11111101011100010011001101100100;
   assign mem[351999:351968] = 32'b11111110000001011010100000111110;
   assign mem[352031:352000] = 32'b00000001001010100100001100001000;
   assign mem[352063:352032] = 32'b00000011011101000001111111001100;
   assign mem[352095:352064] = 32'b11111100000100001011110111011100;
   assign mem[352127:352096] = 32'b11110110000100110011100001110000;
   assign mem[352159:352128] = 32'b00001101000001110011001001000000;
   assign mem[352191:352160] = 32'b11111100100100010100101011010100;
   assign mem[352223:352192] = 32'b00000010010111011110010110111100;
   assign mem[352255:352224] = 32'b11110111001010000000110000110000;
   assign mem[352287:352256] = 32'b11111000110011011111101011101000;
   assign mem[352319:352288] = 32'b00001101000010100111101101110000;
   assign mem[352351:352320] = 32'b11111110011001100100000110000110;
   assign mem[352383:352352] = 32'b11111111110100111001101111001000;
   assign mem[352415:352384] = 32'b11111111000011010101101011010100;
   assign mem[352447:352416] = 32'b00000001000101101010100110100000;
   assign mem[352479:352448] = 32'b00000110010101000101010101101000;
   assign mem[352511:352480] = 32'b11111111100011111100111111000110;
   assign mem[352543:352512] = 32'b00000110010010110000000001110000;
   assign mem[352575:352544] = 32'b11110110010100110101110010000000;
   assign mem[352607:352576] = 32'b11111001100111111110100100010000;
   assign mem[352639:352608] = 32'b11111101111101010111011101111000;
   assign mem[352671:352640] = 32'b00000010100100101101000010000100;
   assign mem[352703:352672] = 32'b11110111000110100100101100000000;
   assign mem[352735:352704] = 32'b00000110011010001101000100000000;
   assign mem[352767:352736] = 32'b11111110110011111100001010001100;
   assign mem[352799:352768] = 32'b00000101000000100110010111100000;
   assign mem[352831:352800] = 32'b11111010101010000010100000010000;
   assign mem[352863:352832] = 32'b00000001011111001000001000101000;
   assign mem[352895:352864] = 32'b11110001001101010010101000100000;
   assign mem[352927:352896] = 32'b00000000010001110110001100001010;
   assign mem[352959:352928] = 32'b00000010101110101010101101101100;
   assign mem[352991:352960] = 32'b11111011011011101100111111100000;
   assign mem[353023:352992] = 32'b00000001011001110000011110010100;
   assign mem[353055:353024] = 32'b00000000010010000110000010001000;
   assign mem[353087:353056] = 32'b11111011000110001010000010000000;
   assign mem[353119:353088] = 32'b11111111110001010110011101111011;
   assign mem[353151:353120] = 32'b11111100101001000101111001001100;
   assign mem[353183:353152] = 32'b11110101000100100000101010110000;
   assign mem[353215:353184] = 32'b11111111110100011001001000111010;
   assign mem[353247:353216] = 32'b00000100001001001111100100001000;
   assign mem[353279:353248] = 32'b00000000110010101100111010011100;
   assign mem[353311:353280] = 32'b11111111011110000110100110100010;
   assign mem[353343:353312] = 32'b11111100100001010101001110000000;
   assign mem[353375:353344] = 32'b00000010101011001110001101011100;
   assign mem[353407:353376] = 32'b00000100011111010011100000100000;
   assign mem[353439:353408] = 32'b11111111100000001110110110011111;
   assign mem[353471:353440] = 32'b00000011100001110110001110011100;
   assign mem[353503:353472] = 32'b00000000110111100011001111000000;
   assign mem[353535:353504] = 32'b11111001001001101101101101011000;
   assign mem[353567:353536] = 32'b00000010000011111011111110001000;
   assign mem[353599:353568] = 32'b00000011010111001000010011101000;
   assign mem[353631:353600] = 32'b11110110110011111001001011110000;
   assign mem[353663:353632] = 32'b00000001010010110111100011110100;
   assign mem[353695:353664] = 32'b11111100011111011100001000101100;
   assign mem[353727:353696] = 32'b11111011111101101110000100110000;
   assign mem[353759:353728] = 32'b00000001101100011100100000000010;
   assign mem[353791:353760] = 32'b11111101100000011111101001001100;
   assign mem[353823:353792] = 32'b00000010010110001100000000010000;
   assign mem[353855:353824] = 32'b00000011110110101110101001000100;
   assign mem[353887:353856] = 32'b11111100011111100100010111000000;
   assign mem[353919:353888] = 32'b00000101101101010010000110111000;
   assign mem[353951:353920] = 32'b11111011011011110010111111011000;
   assign mem[353983:353952] = 32'b00000101110110101101111011010000;
   assign mem[354015:353984] = 32'b11111010111001010111011110011000;
   assign mem[354047:354016] = 32'b00000100001101010101101011111000;
   assign mem[354079:354048] = 32'b00000000100010111100011010010011;
   assign mem[354111:354080] = 32'b00000010010001111000111110010100;
   assign mem[354143:354112] = 32'b00000000110111000100111001000111;
   assign mem[354175:354144] = 32'b11111000000100001100000010111000;
   assign mem[354207:354176] = 32'b11111100000110001001111010011100;
   assign mem[354239:354208] = 32'b00000001001011101111000110110110;
   assign mem[354271:354240] = 32'b00000011011001110100000101101000;
   assign mem[354303:354272] = 32'b11101100110110110011101011100000;
   assign mem[354335:354304] = 32'b00000011010101000011010101011100;
   assign mem[354367:354336] = 32'b00000011100000110010001001101000;
   assign mem[354399:354368] = 32'b00000010001100111110101101010000;
   assign mem[354431:354400] = 32'b11111111000001000000000001010000;
   assign mem[354463:354432] = 32'b00000000000111110001111100101111;
   assign mem[354495:354464] = 32'b11111010001000001010000111110000;
   assign mem[354527:354496] = 32'b11111110000110001010000000101110;
   assign mem[354559:354528] = 32'b00001000000011100011110001100000;
   assign mem[354591:354560] = 32'b11110110001011001000010001000000;
   assign mem[354623:354592] = 32'b00000100101110000101111100011000;
   assign mem[354655:354624] = 32'b11111011110100011000010100001000;
   assign mem[354687:354656] = 32'b11111100001111010110110011101100;
   assign mem[354719:354688] = 32'b11111111011000000001100101110110;
   assign mem[354751:354720] = 32'b11111010110011010010010000111000;
   assign mem[354783:354752] = 32'b11111011100101111011010000001000;
   assign mem[354815:354784] = 32'b00000010010100000001001100111100;
   assign mem[354847:354816] = 32'b00000000001101010000001111010010;
   assign mem[354879:354848] = 32'b00000011110111011100001000101000;
   assign mem[354911:354880] = 32'b00000000111010111101000010011110;
   assign mem[354943:354912] = 32'b11111000110011110010001000111000;
   assign mem[354975:354944] = 32'b11111101110010011000000011111100;
   assign mem[355007:354976] = 32'b11111111100100100011001110010010;
   assign mem[355039:355008] = 32'b11111100010001010000100101010000;
   assign mem[355071:355040] = 32'b11111101110111111001100111100100;
   assign mem[355103:355072] = 32'b11111011110000100110001101111000;
   assign mem[355135:355104] = 32'b00000001110010111011101001000000;
   assign mem[355167:355136] = 32'b11111110100010011001000110011110;
   assign mem[355199:355168] = 32'b00000001001110010110011001100000;
   assign mem[355231:355200] = 32'b00000011001011111001000100110100;
   assign mem[355263:355232] = 32'b11111111100011010000011001010101;
   assign mem[355295:355264] = 32'b00000011001000010011110000100100;
   assign mem[355327:355296] = 32'b11111000000110011010011101111000;
   assign mem[355359:355328] = 32'b11111111011011110011000101000011;
   assign mem[355391:355360] = 32'b11111011000001101110100111111000;
   assign mem[355423:355392] = 32'b11111001100001000010100000010000;
   assign mem[355455:355424] = 32'b11111111010001001011100111100110;
   assign mem[355487:355456] = 32'b00000100101111100110101000110000;
   assign mem[355519:355488] = 32'b00000010000111000001011010111000;
   assign mem[355551:355520] = 32'b00000111100111000111110000000000;
   assign mem[355583:355552] = 32'b00000100110000010110111111110000;
   assign mem[355615:355584] = 32'b11111010001110011110011001111000;
   assign mem[355647:355616] = 32'b00000100111110010001010000010000;
   assign mem[355679:355648] = 32'b11111011010000100100100110010000;
   assign mem[355711:355680] = 32'b11111111111001011011110110001000;
   assign mem[355743:355712] = 32'b00000011000111110101000110101100;
   assign mem[355775:355744] = 32'b11111001011001001010011100010000;
   assign mem[355807:355776] = 32'b00000010110100100100001110111100;
   assign mem[355839:355808] = 32'b11111001111001101001100111100000;
   assign mem[355871:355840] = 32'b00000111111100010101100100010000;
   assign mem[355903:355872] = 32'b00001001100010100110001010000000;
   assign mem[355935:355904] = 32'b11110101011010101011010011000000;
   assign mem[355967:355936] = 32'b00000101000001111100010001101000;
   assign mem[355999:355968] = 32'b11110111000111011101110111100000;
   assign mem[356031:356000] = 32'b00000110011100111011101111100000;
   assign mem[356063:356032] = 32'b00000111010010011001100101110000;
   assign mem[356095:356064] = 32'b11110001001000011001100000000000;
   assign mem[356127:356096] = 32'b00000011101011111100001011001100;
   assign mem[356159:356128] = 32'b11111010010100001100100001011000;
   assign mem[356191:356160] = 32'b00000100111011100101100110000000;
   assign mem[356223:356192] = 32'b00001100110110110001001010100000;
   assign mem[356255:356224] = 32'b00000011000101100110010110101000;
   assign mem[356287:356256] = 32'b11110101110111000110010001110000;
   assign mem[356319:356288] = 32'b11110111100001111010101011010000;
   assign mem[356351:356320] = 32'b11111011100001011010010010011000;
   assign mem[356383:356352] = 32'b11111101100100010100100110100000;
   assign mem[356415:356384] = 32'b00001011101100111100010001110000;
   assign mem[356447:356416] = 32'b11111111110000101101000000001111;
   assign mem[356479:356448] = 32'b11101101100010011001110100100000;
   assign mem[356511:356480] = 32'b00000110110100000001001100111000;
   assign mem[356543:356512] = 32'b11111111001110100011101001011000;
   assign mem[356575:356544] = 32'b00000001000001111001010110101000;
   assign mem[356607:356576] = 32'b11110001101010101011010111100000;
   assign mem[356639:356608] = 32'b00000000010101010000100001001011;
   assign mem[356671:356640] = 32'b00000000110111101010111110001101;
   assign mem[356703:356672] = 32'b00000011110001011100001011110000;
   assign mem[356735:356704] = 32'b11111011111011000101110111101000;
   assign mem[356767:356736] = 32'b00000010110000100111111011010000;
   assign mem[356799:356768] = 32'b11111010001001010011100011010000;
   assign mem[356831:356800] = 32'b00000001110011000100001100010000;
   assign mem[356863:356832] = 32'b00000100000011010001100010110000;
   assign mem[356895:356864] = 32'b00000101001101011011011100110000;
   assign mem[356927:356896] = 32'b11111010110011010110011001110000;
   assign mem[356959:356928] = 32'b11111100000100011110000111110100;
   assign mem[356991:356960] = 32'b11111101100111101010101010001000;
   assign mem[357023:356992] = 32'b11111110101000011001100100010110;
   assign mem[357055:357024] = 32'b00001001101111010010000100000000;
   assign mem[357087:357056] = 32'b11111001110101011111111101011000;
   assign mem[357119:357088] = 32'b11111001001011001000101101010000;
   assign mem[357151:357120] = 32'b00000010001101011100101011010100;
   assign mem[357183:357152] = 32'b11111001000001011111111111100000;
   assign mem[357215:357184] = 32'b00000010110011100110110110101100;
   assign mem[357247:357216] = 32'b11111011110100110001110010100000;
   assign mem[357279:357248] = 32'b00000101111000111110101101001000;
   assign mem[357311:357280] = 32'b11111111001101110010010101010010;
   assign mem[357343:357312] = 32'b11111101101011000000001110100100;
   assign mem[357375:357344] = 32'b11111010000010000111001101000000;
   assign mem[357407:357376] = 32'b00000000010101001000001001101110;
   assign mem[357439:357408] = 32'b00001001000100111010100101000000;
   assign mem[357471:357440] = 32'b00000011111010110100100100111100;
   assign mem[357503:357472] = 32'b00001011101100100000100000100000;
   assign mem[357535:357504] = 32'b00000000010010101010111110100101;
   assign mem[357567:357536] = 32'b00000010000000101011101011010100;
   assign mem[357599:357568] = 32'b00000101000010111100110110101000;
   assign mem[357631:357600] = 32'b00000000000110100001110101110010;
   assign mem[357663:357632] = 32'b11111110000110010101111011100110;
   assign mem[357695:357664] = 32'b00001000110010111000101011000000;
   assign mem[357727:357696] = 32'b11110010111000111011100110100000;
   assign mem[357759:357728] = 32'b11111100011011110101011011000000;
   assign mem[357791:357760] = 32'b00000101000000100001000011000000;
   assign mem[357823:357792] = 32'b00000011010000001110010110011000;
   assign mem[357855:357824] = 32'b11111111010011011010010000110111;
   assign mem[357887:357856] = 32'b11110111100111110100011110000000;
   assign mem[357919:357888] = 32'b11111111000110101100101111110101;
   assign mem[357951:357920] = 32'b11111111101110010110111101001000;
   assign mem[357983:357952] = 32'b00000101110111100001011001000000;
   assign mem[358015:357984] = 32'b11111110000111101110011101001000;
   assign mem[358047:358016] = 32'b00000000110111001011110011011010;
   assign mem[358079:358048] = 32'b00000000001011101010000101001111;
   assign mem[358111:358080] = 32'b11111100110111111000100000011100;
   assign mem[358143:358112] = 32'b11111001111000001110101010101000;
   assign mem[358175:358144] = 32'b11111111010101001011101111000100;
   assign mem[358207:358176] = 32'b00000010110110000011010010001100;
   assign mem[358239:358208] = 32'b00000100100101101101100100111000;
   assign mem[358271:358240] = 32'b00000001011001011100101000000100;
   assign mem[358303:358272] = 32'b00000001010011001110000111101010;
   assign mem[358335:358304] = 32'b11111111001001010101100101010110;
   assign mem[358367:358336] = 32'b11111011000101000111111111011000;
   assign mem[358399:358368] = 32'b00000100001111110001000100110000;
   assign mem[358431:358400] = 32'b11111001010111100110000100011000;
   assign mem[358463:358432] = 32'b11111110000001101101111000111010;
   assign mem[358495:358464] = 32'b00000100000001000011011000011000;
   assign mem[358527:358496] = 32'b11111111101000110010110100010001;
   assign mem[358559:358528] = 32'b11111001100100011001010101100000;
   assign mem[358591:358560] = 32'b11111110001010100100010101010100;
   assign mem[358623:358592] = 32'b00000010001001011110001111111100;
   assign mem[358655:358624] = 32'b00000010100111011100100001001000;
   assign mem[358687:358656] = 32'b00000011011000100111101111001100;
   assign mem[358719:358688] = 32'b11111111001011101010001101011101;
   assign mem[358751:358720] = 32'b11111111100111101010010000011010;
   assign mem[358783:358752] = 32'b00000101100000111011011010101000;
   assign mem[358815:358784] = 32'b00000101001110010110010010111000;
   assign mem[358847:358816] = 32'b11111011000000100100000101011000;
   assign mem[358879:358848] = 32'b00000010011010000011011011011100;
   assign mem[358911:358880] = 32'b00000100100111111101111101111000;
   assign mem[358943:358912] = 32'b11111111110010111011000001011011;
   assign mem[358975:358944] = 32'b00000010001100010010011100110000;
   assign mem[359007:358976] = 32'b11111001010100111101111110101000;
   assign mem[359039:359008] = 32'b11111111010101101011100000110001;
   assign mem[359071:359040] = 32'b11111010000010110100110011010000;
   assign mem[359103:359072] = 32'b11111101000000011010110001110100;
   assign mem[359135:359104] = 32'b00000000101110000111000000110100;
   assign mem[359167:359136] = 32'b00000000110001001110100001110101;
   assign mem[359199:359168] = 32'b00000110011011100101101101110000;
   assign mem[359231:359200] = 32'b00000000000111011101111000110100;
   assign mem[359263:359232] = 32'b11111111100100100001100110000101;
   assign mem[359295:359264] = 32'b11111011110101010111100111000000;
   assign mem[359327:359296] = 32'b11111110001110101011000000101010;
   assign mem[359359:359328] = 32'b00000000001000111010100111101001;
   assign mem[359391:359360] = 32'b00001010100001111001110011110000;
   assign mem[359423:359392] = 32'b00011000001110101100011010100000;
   assign mem[359455:359424] = 32'b00000010000110011110111101001000;
   assign mem[359487:359456] = 32'b11111100010010011100110000010100;
   assign mem[359519:359488] = 32'b11110001001110110000001110010000;
   assign mem[359551:359520] = 32'b11111110101110010011101101101110;
   assign mem[359583:359552] = 32'b11111101111001111111111100011100;
   assign mem[359615:359584] = 32'b00001110011010011000010010000000;
   assign mem[359647:359616] = 32'b11111000110010011011100010010000;
   assign mem[359679:359648] = 32'b11101111111101111010101111100000;
   assign mem[359711:359680] = 32'b00000100110110111010001110000000;
   assign mem[359743:359712] = 32'b11111010100100110100101110011000;
   assign mem[359775:359744] = 32'b11111011100001011101101011001000;
   assign mem[359807:359776] = 32'b00001000010000001001100001100000;
   assign mem[359839:359808] = 32'b11111111011110011100001001010101;
   assign mem[359871:359840] = 32'b00000010110100010110001001010000;
   assign mem[359903:359872] = 32'b11111010010010111010011101101000;
   assign mem[359935:359904] = 32'b11111000110010001011010000000000;
   assign mem[359967:359936] = 32'b11111101110011001000110000000100;
   assign mem[359999:359968] = 32'b00000010101000111000000110011100;
   assign mem[360031:360000] = 32'b00000011101001000111111110011000;
   assign mem[360063:360032] = 32'b11110010100110000110100001100000;
   assign mem[360095:360064] = 32'b00000010001010001011100110110000;
   assign mem[360127:360096] = 32'b11111101000111111011000001110100;
   assign mem[360159:360128] = 32'b11111111101011000011111010011110;
   assign mem[360191:360160] = 32'b00000110111011101100100101110000;
   assign mem[360223:360192] = 32'b00000011011000011101010011100000;
   assign mem[360255:360224] = 32'b11110111101001011010101100010000;
   assign mem[360287:360256] = 32'b11111001011111011111101011001000;
   assign mem[360319:360288] = 32'b00000001011111010110001100100000;
   assign mem[360351:360320] = 32'b11111110000001001000101111000100;
   assign mem[360383:360352] = 32'b11110111101011011000001001110000;
   assign mem[360415:360384] = 32'b00000010001010001101100000100000;
   assign mem[360447:360416] = 32'b11111100111011010101011010100100;
   assign mem[360479:360448] = 32'b00000101101100011000000011010000;
   assign mem[360511:360480] = 32'b00000010001111001100011010000100;
   assign mem[360543:360512] = 32'b11111111101000111000101001000010;
   assign mem[360575:360544] = 32'b11110001110101101000000000010000;
   assign mem[360607:360576] = 32'b11111110011101011101111011100110;
   assign mem[360639:360608] = 32'b00000110110000000110011011011000;
   assign mem[360671:360640] = 32'b11111010100010101110100110011000;
   assign mem[360703:360672] = 32'b11110100100101110101100001000000;
   assign mem[360735:360704] = 32'b11110101111011100010011111110000;
   assign mem[360767:360736] = 32'b00000111110101100011011000100000;
   assign mem[360799:360768] = 32'b00000100011001111101000100101000;
   assign mem[360831:360800] = 32'b00000001111100111111100110110110;
   assign mem[360863:360832] = 32'b11110101000110000011010010000000;
   assign mem[360895:360864] = 32'b00000001101110110010011111000010;
   assign mem[360927:360896] = 32'b11111010010101010110111001100000;
   assign mem[360959:360928] = 32'b00001000100000010111111000010000;
   assign mem[360991:360960] = 32'b11110100011110110101101011110000;
   assign mem[361023:360992] = 32'b00000111101000110111100110100000;
   assign mem[361055:361024] = 32'b00000100000001001101001100010000;
   assign mem[361087:361056] = 32'b00000110001100111000011001000000;
   assign mem[361119:361088] = 32'b00000000011000101101001111010101;
   assign mem[361151:361120] = 32'b00000001000111100101000110111010;
   assign mem[361183:361152] = 32'b11111100010011101110100000011000;
   assign mem[361215:361184] = 32'b11111000011001101000101110011000;
   assign mem[361247:361216] = 32'b00000000100111001110100000101111;
   assign mem[361279:361248] = 32'b11111101110001010101010010000100;
   assign mem[361311:361280] = 32'b11101100101001100101010010100000;
   assign mem[361343:361312] = 32'b00000110101000101100001101000000;
   assign mem[361375:361344] = 32'b00000001010100000110101111001000;
   assign mem[361407:361376] = 32'b00000011101011100100001011001100;
   assign mem[361439:361408] = 32'b00000010100100001010111010110000;
   assign mem[361471:361440] = 32'b00000011100111100111100011100100;
   assign mem[361503:361472] = 32'b11111010101111110000010111111000;
   assign mem[361535:361504] = 32'b11111011010101010100010101001000;
   assign mem[361567:361536] = 32'b11111110010111001011100101001000;
   assign mem[361599:361568] = 32'b00000101001100000111000110000000;
   assign mem[361631:361600] = 32'b11111000000000111100110100111000;
   assign mem[361663:361632] = 32'b11110100111110000000110100000000;
   assign mem[361695:361664] = 32'b11111001101101100001001101001000;
   assign mem[361727:361696] = 32'b00001011001110111111010000010000;
   assign mem[361759:361728] = 32'b00000100000101001000000110110000;
   assign mem[361791:361760] = 32'b00000001110100011100100110011110;
   assign mem[361823:361792] = 32'b11111011000110110000111110000000;
   assign mem[361855:361824] = 32'b11111000111011000110110000100000;
   assign mem[361887:361856] = 32'b11110110110010010110111000000000;
   assign mem[361919:361888] = 32'b00000110100010011101111001111000;
   assign mem[361951:361920] = 32'b00001000110111000100011010100000;
   assign mem[361983:361952] = 32'b00000010001011000111010111110000;
   assign mem[362015:361984] = 32'b00000001100100001110111011000010;
   assign mem[362047:362016] = 32'b00000011100001101010101000110000;
   assign mem[362079:362048] = 32'b11110111111101111110001000110000;
   assign mem[362111:362080] = 32'b00000000111100000010001001011001;
   assign mem[362143:362112] = 32'b00000110000110000001011011111000;
   assign mem[362175:362144] = 32'b11111011010010110001011000001000;
   assign mem[362207:362176] = 32'b00000111100001110001100000001000;
   assign mem[362239:362208] = 32'b11101111111011110101111101000000;
   assign mem[362271:362240] = 32'b11111100100111010010110010001000;
   assign mem[362303:362272] = 32'b11111100011001001101001101011000;
   assign mem[362335:362304] = 32'b00000011101011000111110111110100;
   assign mem[362367:362336] = 32'b00000011101110110010001111001000;
   assign mem[362399:362368] = 32'b00000111010101001010111100011000;
   assign mem[362431:362400] = 32'b11111111101001110010100111100110;
   assign mem[362463:362432] = 32'b00001001110101010111110010110000;
   assign mem[362495:362464] = 32'b11111011011111110101100011101000;
   assign mem[362527:362496] = 32'b11111000101110110010011011100000;
   assign mem[362559:362528] = 32'b11111110001010100110110111010100;
   assign mem[362591:362560] = 32'b11110100010100010111011010110000;
   assign mem[362623:362592] = 32'b00000011001000000101010010110000;
   assign mem[362655:362624] = 32'b11111110110001001100111010000010;
   assign mem[362687:362656] = 32'b11111101110110101010101110010000;
   assign mem[362719:362688] = 32'b00000011110011010001000011100000;
   assign mem[362751:362720] = 32'b00000101011101000011011011101000;
   assign mem[362783:362752] = 32'b00000000111011101101101110010100;
   assign mem[362815:362784] = 32'b11111010111100111100001010101000;
   assign mem[362847:362816] = 32'b00000110010010100101110010011000;
   assign mem[362879:362848] = 32'b11111010010010011011110010011000;
   assign mem[362911:362880] = 32'b11101010010100111101101000100000;
   assign mem[362943:362912] = 32'b00001100100100000110101011110000;
   assign mem[362975:362944] = 32'b11111100010000110100101000000000;
   assign mem[363007:362976] = 32'b11111011101011111101101100010000;
   assign mem[363039:363008] = 32'b00001000011100010110100000010000;
   assign mem[363071:363040] = 32'b11111111010000110000000100111110;
   assign mem[363103:363072] = 32'b11110111110101111011010101110000;
   assign mem[363135:363104] = 32'b00000001001101000010011010111000;
   assign mem[363167:363136] = 32'b11111101100101100110111111000100;
   assign mem[363199:363168] = 32'b00000011101111101001011001101100;
   assign mem[363231:363200] = 32'b11111100110111111001010001011000;
   assign mem[363263:363232] = 32'b00000001100001100101011001100110;
   assign mem[363295:363264] = 32'b11111111101110001000100011110111;
   assign mem[363327:363296] = 32'b11111111101100011000001010011110;
   assign mem[363359:363328] = 32'b11111101101111011011011010011100;
   assign mem[363391:363360] = 32'b11111111101101111111011100010110;
   assign mem[363423:363392] = 32'b00000001100110100110010000100110;
   assign mem[363455:363424] = 32'b00000000010011100111001010011011;
   assign mem[363487:363456] = 32'b11111011111000111011010010010000;
   assign mem[363519:363488] = 32'b00000010011001011000101010101000;
   assign mem[363551:363520] = 32'b11110011010010110110100001110000;
   assign mem[363583:363552] = 32'b00000100110110101000101001110000;
   assign mem[363615:363584] = 32'b00000101010100100011001000100000;
   assign mem[363647:363616] = 32'b11111011101100010101001110000000;
   assign mem[363679:363648] = 32'b11111010011011100100011000111000;
   assign mem[363711:363680] = 32'b11111011000001100000111011110000;
   assign mem[363743:363712] = 32'b00000000001100000011010011101001;
   assign mem[363775:363744] = 32'b00000101011110010111010000001000;
   assign mem[363807:363776] = 32'b00000011111101101111111011011100;
   assign mem[363839:363808] = 32'b11110100011001010100111010000000;
   assign mem[363871:363840] = 32'b11111100010100101010010001000100;
   assign mem[363903:363872] = 32'b00000010000111001001000010000100;
   assign mem[363935:363904] = 32'b00000010011110110011110001010100;
   assign mem[363967:363936] = 32'b11111110101000001101010011101100;
   assign mem[363999:363968] = 32'b00000001101010010011000000000000;
   assign mem[364031:364000] = 32'b11111101011111110101101101111100;
   assign mem[364063:364032] = 32'b00000000100111001000011110110111;
   assign mem[364095:364064] = 32'b11111111000000000110111111111101;
   assign mem[364127:364096] = 32'b11111101010000101110001100011100;
   assign mem[364159:364128] = 32'b11111101111110011111101001001000;
   assign mem[364191:364160] = 32'b00001000011011011110100110000000;
   assign mem[364223:364192] = 32'b11111000000011010100010110111000;
   assign mem[364255:364224] = 32'b00000010100110010101000000100000;
   assign mem[364287:364256] = 32'b11111101000011010111100100110100;
   assign mem[364319:364288] = 32'b00000000110000101010001101011110;
   assign mem[364351:364320] = 32'b11111100011111110111000111010100;
   assign mem[364383:364352] = 32'b00000000010100110000011111110100;
   assign mem[364415:364384] = 32'b11111111001101101011000110011010;
   assign mem[364447:364416] = 32'b00000001001000001010001010001010;
   assign mem[364479:364448] = 32'b00000011001100001011111100101000;
   assign mem[364511:364480] = 32'b11110000001011011110111110110000;
   assign mem[364543:364512] = 32'b00001011111100101111110111010000;
   assign mem[364575:364544] = 32'b11110100100100001111111011110000;
   assign mem[364607:364576] = 32'b00000101001001110111101101110000;
   assign mem[364639:364608] = 32'b00000010011010000000000100000000;
   assign mem[364671:364640] = 32'b00000011010011010010010110010000;
   assign mem[364703:364672] = 32'b11111010111101110110000000001000;
   assign mem[364735:364704] = 32'b00000011011110100010110110100000;
   assign mem[364767:364736] = 32'b11110001011000110000000100100000;
   assign mem[364799:364768] = 32'b00000100101011101000001110001000;
   assign mem[364831:364800] = 32'b11111101010001001011101001101100;
   assign mem[364863:364832] = 32'b11110110010000101011000001010000;
   assign mem[364895:364864] = 32'b11111010111010001001110011010000;
   assign mem[364927:364896] = 32'b00000000111001111000100011110110;
   assign mem[364959:364928] = 32'b00000010011100100101101000101100;
   assign mem[364991:364960] = 32'b11111100111011101110001000110100;
   assign mem[365023:364992] = 32'b11111110001100101000000110001010;
   assign mem[365055:365024] = 32'b00000000101111101011010111010110;
   assign mem[365087:365056] = 32'b11111101011000111011010110111100;
   assign mem[365119:365088] = 32'b00000100100011111100010111110000;
   assign mem[365151:365120] = 32'b11111110010100101000010001101000;
   assign mem[365183:365152] = 32'b11110100110001001001100110100000;
   assign mem[365215:365184] = 32'b11111110010100011011111111101110;
   assign mem[365247:365216] = 32'b00000100011011100110101001010000;
   assign mem[365279:365248] = 32'b00000100111000100011001100000000;
   assign mem[365311:365280] = 32'b00000000011010111001011010110000;
   assign mem[365343:365312] = 32'b11111111000011101110000000011101;
   assign mem[365375:365344] = 32'b11111111110111001110000101101010;
   assign mem[365407:365376] = 32'b11111000101011000100100110111000;
   assign mem[365439:365408] = 32'b11111110110010001010101101001110;
   assign mem[365471:365440] = 32'b00000000100100001100001011001100;
   assign mem[365503:365472] = 32'b00000001010011101011111000010010;
   assign mem[365535:365504] = 32'b00000010110111111110101010000100;
   assign mem[365567:365536] = 32'b00000111111001101110101001110000;
   assign mem[365599:365568] = 32'b11111011110100101001110111001000;
   assign mem[365631:365600] = 32'b11111011011100000100011111110000;
   assign mem[365663:365632] = 32'b00000000000010100000000110011111;
   assign mem[365695:365664] = 32'b11111101111010011101100010100000;
   assign mem[365727:365696] = 32'b11111111100101010000000101001001;
   assign mem[365759:365728] = 32'b11111100011110000100111011111100;
   assign mem[365791:365760] = 32'b00001111100010011111110111010000;
   assign mem[365823:365792] = 32'b00000001110011010111101001110100;
   assign mem[365855:365824] = 32'b11111111010001101011101011001001;
   assign mem[365887:365856] = 32'b11101110111110010101011111000000;
   assign mem[365919:365888] = 32'b11111001000101101111001000100000;
   assign mem[365951:365920] = 32'b00000000001111001101010010110100;
   assign mem[365983:365952] = 32'b11111101010011111010110011001000;
   assign mem[366015:365984] = 32'b00000000101001010110111010010111;
   assign mem[366047:366016] = 32'b00000011010010000100010101000000;
   assign mem[366079:366048] = 32'b11111001010011001101010011111000;
   assign mem[366111:366080] = 32'b00000000110110111101001100011010;
   assign mem[366143:366112] = 32'b00001100000101101000001101100000;
   assign mem[366175:366144] = 32'b11111011110010011101011001001000;
   assign mem[366207:366176] = 32'b00000110001001110010010100010000;
   assign mem[366239:366208] = 32'b00000000111111011111110110101101;
   assign mem[366271:366240] = 32'b00000001001011100001101111011000;
   assign mem[366303:366272] = 32'b00000100101101010100100110001000;
   assign mem[366335:366304] = 32'b11111011010110001011000010000000;
   assign mem[366367:366336] = 32'b11111101011010110110111010100100;
   assign mem[366399:366368] = 32'b11110100001100101110101011000000;
   assign mem[366431:366400] = 32'b11110001001001000001011010110000;
   assign mem[366463:366432] = 32'b11111010010110111010011110010000;
   assign mem[366495:366464] = 32'b11111110110011110010011100011110;
   assign mem[366527:366496] = 32'b00000000001101010111011111000101;
   assign mem[366559:366528] = 32'b00001000101001111010111010000000;
   assign mem[366591:366560] = 32'b00000011100000001100110110110000;
   assign mem[366623:366592] = 32'b11111000011111001001111000001000;
   assign mem[366655:366624] = 32'b11111010110011111000100000001000;
   assign mem[366687:366656] = 32'b11111111100100110101001110101101;
   assign mem[366719:366688] = 32'b00000011001100111100111011110100;
   assign mem[366751:366720] = 32'b00000101100101100111100110110000;
   assign mem[366783:366752] = 32'b00000010101011000111011011101000;
   assign mem[366815:366784] = 32'b00000010010011000110100011010100;
   assign mem[366847:366816] = 32'b00000101101000001101011110001000;
   assign mem[366879:366848] = 32'b11111101000011010111110000100100;
   assign mem[366911:366880] = 32'b00000001000110001000010100100110;
   assign mem[366943:366912] = 32'b11111010110000011101110101110000;
   assign mem[366975:366944] = 32'b11111010111011100010111000101000;
   assign mem[367007:366976] = 32'b11110000010000001111001110110000;
   assign mem[367039:367008] = 32'b11111110101100101011101110110000;
   assign mem[367071:367040] = 32'b11111101000011111110000000100100;
   assign mem[367103:367072] = 32'b00000100101111011010101100011000;
   assign mem[367135:367104] = 32'b00000001010010011000010111111100;
   assign mem[367167:367136] = 32'b00000011001000011110011100000100;
   assign mem[367199:367168] = 32'b11111011010110101011100000000000;
   assign mem[367231:367200] = 32'b00000010101011101001000110000100;
   assign mem[367263:367232] = 32'b00001000010010011101011011010000;
   assign mem[367295:367264] = 32'b11111010011101101101011010101000;
   assign mem[367327:367296] = 32'b00001001000111101011111000100000;
   assign mem[367359:367328] = 32'b11110110010111010110010100110000;
   assign mem[367391:367360] = 32'b00000011010101001001111001101000;
   assign mem[367423:367392] = 32'b11111100000101110101010011001000;
   assign mem[367455:367424] = 32'b00000101100101111000110000111000;
   assign mem[367487:367456] = 32'b11111111110100101001010110001110;
   assign mem[367519:367488] = 32'b11111011000001010111010011111000;
   assign mem[367551:367520] = 32'b00000011110011000010001111010100;
   assign mem[367583:367552] = 32'b11110110000111000100000100010000;
   assign mem[367615:367584] = 32'b00000101010011101001001110001000;
   assign mem[367647:367616] = 32'b11111000110100000101001110011000;
   assign mem[367679:367648] = 32'b00000001001111111110110000010100;
   assign mem[367711:367680] = 32'b11111111011101101011010100110010;
   assign mem[367743:367712] = 32'b00000010000101011001111011100000;
   assign mem[367775:367744] = 32'b00000101100000010100010011101000;
   assign mem[367807:367776] = 32'b11111110001011010111110010000100;
   assign mem[367839:367808] = 32'b11111100100001111101000101111100;
   assign mem[367871:367840] = 32'b00000000111001011000101111100000;
   assign mem[367903:367872] = 32'b00000011001111100100111100011100;
   assign mem[367935:367904] = 32'b00000000100010001110000010101000;
   assign mem[367967:367936] = 32'b11111111100110001001101100100100;
   assign mem[367999:367968] = 32'b00000011111010110001011011010000;
   assign mem[368031:368000] = 32'b11110101111011011110001001010000;
   assign mem[368063:368032] = 32'b00000111101011101000110100111000;
   assign mem[368095:368064] = 32'b11111001110011110010000011011000;
   assign mem[368127:368096] = 32'b00000001010101110010010110111010;
   assign mem[368159:368128] = 32'b11110111110101000011000010100000;
   assign mem[368191:368160] = 32'b00000001111111010010100010001010;
   assign mem[368223:368192] = 32'b11111111110111111110111111000001;
   assign mem[368255:368224] = 32'b00000010011111111001101111100000;
   assign mem[368287:368256] = 32'b11111001101111000001111100010000;
   assign mem[368319:368288] = 32'b11111111101010001100111000011001;
   assign mem[368351:368320] = 32'b11111100100000010110000100011100;
   assign mem[368383:368352] = 32'b00000111010011101011111010101000;
   assign mem[368415:368384] = 32'b00000101000111100101110100001000;
   assign mem[368447:368416] = 32'b11111101110000111001001001001000;
   assign mem[368479:368448] = 32'b11111110101101100101110110101000;
   assign mem[368511:368480] = 32'b11111111010011111111000000010011;
   assign mem[368543:368512] = 32'b00000100001101101000111100011000;
   assign mem[368575:368544] = 32'b11111111100000110010111110000010;
   assign mem[368607:368576] = 32'b11111011101101000001001101001000;
   assign mem[368639:368608] = 32'b11111110010111011010100101101000;
   assign mem[368671:368640] = 32'b00000010001010000011001101011100;
   assign mem[368703:368672] = 32'b11110110011110001101010011100000;
   assign mem[368735:368704] = 32'b00000010010000101000000101110100;
   assign mem[368767:368736] = 32'b11111111100101000001001011100010;
   assign mem[368799:368768] = 32'b11111101010000101000110011111000;
   assign mem[368831:368800] = 32'b00000000010000001101000111001111;
   assign mem[368863:368832] = 32'b00000000101001011011011011011111;
   assign mem[368895:368864] = 32'b00000001101100000001110001110110;
   assign mem[368927:368896] = 32'b00000111010011001101011010110000;
   assign mem[368959:368928] = 32'b11111000101000011000101100111000;
   assign mem[368991:368960] = 32'b11111100100111111010010111011100;
   assign mem[369023:368992] = 32'b00000001111001010101100000111100;
   assign mem[369055:369024] = 32'b11110100101100101110101100110000;
   assign mem[369087:369056] = 32'b00000011111101100110010110001000;
   assign mem[369119:369088] = 32'b11101000010010011010000101000000;
   assign mem[369151:369120] = 32'b00000111111001111000000011111000;
   assign mem[369183:369152] = 32'b00001100111001100101001011000000;
   assign mem[369215:369184] = 32'b11110000100111111100011000100000;
   assign mem[369247:369216] = 32'b00000010000000010001000000111100;
   assign mem[369279:369248] = 32'b11111001011001111001011100110000;
   assign mem[369311:369280] = 32'b11110111100011010101001000110000;
   assign mem[369343:369312] = 32'b11111110010011110001110010010100;
   assign mem[369375:369344] = 32'b00000101011110000110000011011000;
   assign mem[369407:369376] = 32'b00000110110100110000000101011000;
   assign mem[369439:369408] = 32'b11111001011000100000100100111000;
   assign mem[369471:369440] = 32'b00000111011001010010100100011000;
   assign mem[369503:369472] = 32'b00000001001010110010010110101110;
   assign mem[369535:369504] = 32'b11110101000001000110011111000000;
   assign mem[369567:369536] = 32'b00000010001100000101111110111000;
   assign mem[369599:369568] = 32'b11110101000111101110011111100000;
   assign mem[369631:369600] = 32'b11111110000001010111111011010100;
   assign mem[369663:369632] = 32'b11110011000101011100000001000000;
   assign mem[369695:369664] = 32'b00000000100111001011111010001110;
   assign mem[369727:369696] = 32'b00000011111101111101110111110100;
   assign mem[369759:369728] = 32'b11111101101011000110100101111000;
   assign mem[369791:369760] = 32'b11111111010000100010000001010000;
   assign mem[369823:369792] = 32'b11111110110111001111010111010000;
   assign mem[369855:369824] = 32'b11111100000101000101000101011000;
   assign mem[369887:369856] = 32'b11111101011001110111011011001100;
   assign mem[369919:369888] = 32'b11111110001101001011111000011000;
   assign mem[369951:369920] = 32'b00000000101101010001000001101010;
   assign mem[369983:369952] = 32'b00001000111011011101001001010000;
   assign mem[370015:369984] = 32'b11111101010111001101100110111100;
   assign mem[370047:370016] = 32'b00000000010001110100111000010001;
   assign mem[370079:370048] = 32'b11111101101011111011010011111000;
   assign mem[370111:370080] = 32'b11110111101110100011000100110000;
   assign mem[370143:370112] = 32'b11110111001010011000101100110000;
   assign mem[370175:370144] = 32'b00000010110100001000010011001100;
   assign mem[370207:370176] = 32'b00000101111110111001000011001000;
   assign mem[370239:370208] = 32'b11111110100101011010110011111010;
   assign mem[370271:370240] = 32'b11111111101001010011111111000100;
   assign mem[370303:370272] = 32'b00000001111110110000101000100100;
   assign mem[370335:370304] = 32'b00000010101001001100100111010100;
   assign mem[370367:370336] = 32'b11111101010110001001100011010000;
   assign mem[370399:370368] = 32'b11111011111010011110011001100000;
   assign mem[370431:370400] = 32'b00000010000011011001000010011000;
   assign mem[370463:370432] = 32'b00000001010000000100101010100110;
   assign mem[370495:370464] = 32'b00000100010001011011110010111000;
   assign mem[370527:370496] = 32'b11111000011000011000000111001000;
   assign mem[370559:370528] = 32'b11111111011110000100100011011000;
   assign mem[370591:370560] = 32'b11111010111010111011100011011000;
   assign mem[370623:370592] = 32'b00000100111101111000111010110000;
   assign mem[370655:370624] = 32'b11111110011101010101100000011100;
   assign mem[370687:370656] = 32'b00000001111011100110011110001010;
   assign mem[370719:370688] = 32'b11111011111110101000010101011000;
   assign mem[370751:370720] = 32'b00000001011010001101001101011110;
   assign mem[370783:370752] = 32'b11111010111101011000000011101000;
   assign mem[370815:370784] = 32'b11111111100010000100100111000101;
   assign mem[370847:370816] = 32'b11111110101010011011111111001000;
   assign mem[370879:370848] = 32'b00000001100001011000110011000010;
   assign mem[370911:370880] = 32'b00000101111100011010001111010000;
   assign mem[370943:370912] = 32'b11111010100010010100101001101000;
   assign mem[370975:370944] = 32'b00000001001101011110011000000000;
   assign mem[371007:370976] = 32'b00000011010001010001101010010000;
   assign mem[371039:371008] = 32'b11111011011101100010000101110000;
   assign mem[371071:371040] = 32'b11111100010001110101010000011000;
   assign mem[371103:371072] = 32'b00000000110010110011000011111101;
   assign mem[371135:371104] = 32'b00000000111101001011001010010001;
   assign mem[371167:371136] = 32'b00000100101000011111111110110000;
   assign mem[371199:371168] = 32'b00000000101111111100100001001011;
   assign mem[371231:371200] = 32'b00010000101000000111011011100000;
   assign mem[371263:371232] = 32'b11110010001110010101000111110000;
   assign mem[371295:371264] = 32'b00000010011110010100101010011000;
   assign mem[371327:371296] = 32'b11111100010011101000100000101000;
   assign mem[371359:371328] = 32'b11110100011011000001000100010000;
   assign mem[371391:371360] = 32'b00000010011001100111100111101000;
   assign mem[371423:371392] = 32'b00000010010101010011101111101100;
   assign mem[371455:371424] = 32'b00000101110010000001011001110000;
   assign mem[371487:371456] = 32'b11111001011110101010000111101000;
   assign mem[371519:371488] = 32'b11110000000101110011100101010000;
   assign mem[371551:371520] = 32'b00000001000111100011010110000010;
   assign mem[371583:371552] = 32'b00010110100101011000001000100000;
   assign mem[371615:371584] = 32'b11110101011100000110100011100000;
   assign mem[371647:371616] = 32'b00000001000110011010010100010010;
   assign mem[371679:371648] = 32'b11111111101010110111101100101001;
   assign mem[371711:371680] = 32'b00001000110111010101011000110000;
   assign mem[371743:371712] = 32'b11110110011010010011011000000000;
   assign mem[371775:371744] = 32'b00001000001010110111101011100000;
   assign mem[371807:371776] = 32'b11110101011000011011111011010000;
   assign mem[371839:371808] = 32'b11111101010100111001101101000100;
   assign mem[371871:371840] = 32'b00000011001001111100000010011000;
   assign mem[371903:371872] = 32'b11111010100000000110110100000000;
   assign mem[371935:371904] = 32'b00000001000101100110010100100110;
   assign mem[371967:371936] = 32'b11111000010100011000010110101000;
   assign mem[371999:371968] = 32'b00000001100010010111111001010000;
   assign mem[372031:372000] = 32'b11111110001010110011100010001100;
   assign mem[372063:372032] = 32'b00000000100011001110000101111101;
   assign mem[372095:372064] = 32'b00000010000011110111000011101100;
   assign mem[372127:372096] = 32'b00001001001011101111001111110000;
   assign mem[372159:372128] = 32'b00000100110010110011010110010000;
   assign mem[372191:372160] = 32'b00000001010110000001000110110010;
   assign mem[372223:372192] = 32'b11111100001001101100000111101100;
   assign mem[372255:372224] = 32'b11111110001110111001000110010000;
   assign mem[372287:372256] = 32'b00000101101010010010011110101000;
   assign mem[372319:372288] = 32'b11111101100110110000011010010100;
   assign mem[372351:372320] = 32'b00000110001000100000101100110000;
   assign mem[372383:372352] = 32'b00000001010000011110011100110110;
   assign mem[372415:372384] = 32'b11111011000010011101011101000000;
   assign mem[372447:372416] = 32'b00000010000101010111100111011000;
   assign mem[372479:372448] = 32'b11111111000111000001111110111100;
   assign mem[372511:372480] = 32'b11111110001100101111011101111110;
   assign mem[372543:372512] = 32'b00000100100001101011110101001000;
   assign mem[372575:372544] = 32'b00001000010000100011100111010000;
   assign mem[372607:372576] = 32'b11111011001011111101110011000000;
   assign mem[372639:372608] = 32'b00001000000010100100110100000000;
   assign mem[372671:372640] = 32'b11110111001101010000001100010000;
   assign mem[372703:372672] = 32'b00000000000110000110101110111101;
   assign mem[372735:372704] = 32'b00000100110011110000101100000000;
   assign mem[372767:372736] = 32'b11110111100010110100010000000000;
   assign mem[372799:372768] = 32'b11111001101100110000010110100000;
   assign mem[372831:372800] = 32'b00000101101000100101000100110000;
   assign mem[372863:372832] = 32'b11111010001011110110011001011000;
   assign mem[372895:372864] = 32'b00000110011111010110111000101000;
   assign mem[372927:372896] = 32'b00000110111001100010011100001000;
   assign mem[372959:372928] = 32'b11110011111110100111110100100000;
   assign mem[372991:372960] = 32'b00000011000000001110100010100000;
   assign mem[373023:372992] = 32'b00000100010101101110000000011000;
   assign mem[373055:373024] = 32'b00000000100001000000101000010110;
   assign mem[373087:373056] = 32'b00000000001110110111111111011000;
   assign mem[373119:373088] = 32'b11100100100000110111011111100000;
   assign mem[373151:373120] = 32'b11110011011110000101101001110000;
   assign mem[373183:373152] = 32'b00000100010001110001110101111000;
   assign mem[373215:373184] = 32'b00000011101011101111110110110100;
   assign mem[373247:373216] = 32'b00000010000100011111010001101000;
   assign mem[373279:373248] = 32'b00000001010011000001101111000000;
   assign mem[373311:373280] = 32'b11111011100010001011111100010000;
   assign mem[373343:373312] = 32'b00000100010010001100001101000000;
   assign mem[373375:373344] = 32'b11111110000010011101000001000000;
   assign mem[373407:373376] = 32'b00000110101100111110001010101000;
   assign mem[373439:373408] = 32'b11110111110110010110100111000000;
   assign mem[373471:373440] = 32'b00000001000000010000010111010100;
   assign mem[373503:373472] = 32'b11110100010101001100000000110000;
   assign mem[373535:373504] = 32'b00000010001001001110010101101100;
   assign mem[373567:373536] = 32'b00000010111000110000100110111100;
   assign mem[373599:373568] = 32'b11111010100001101101100111100000;
   assign mem[373631:373600] = 32'b00000100000010111001101111001000;
   assign mem[373663:373632] = 32'b11111111111000101100101110010101;
   assign mem[373695:373664] = 32'b00000000101100111101100010100000;
   assign mem[373727:373696] = 32'b00000000000010000101100101011010;
   assign mem[373759:373728] = 32'b11111011000001000100010000011000;
   assign mem[373791:373760] = 32'b00000010101010111110001111010100;
   assign mem[373823:373792] = 32'b00000011101011111000110111000100;
   assign mem[373855:373824] = 32'b11111001010010100111100111010000;
   assign mem[373887:373856] = 32'b11111100001011011111010011111000;
   assign mem[373919:373888] = 32'b00000100110011101011011100110000;
   assign mem[373951:373920] = 32'b11110110011111101101010101110000;
   assign mem[373983:373952] = 32'b00001001111111110011000010110000;
   assign mem[374015:373984] = 32'b11111111110011111111100100101111;
   assign mem[374047:374016] = 32'b11111101010011000010110001110000;
   assign mem[374079:374048] = 32'b00000011001001100100001101110000;
   assign mem[374111:374080] = 32'b11110101100101001000011010010000;
   assign mem[374143:374112] = 32'b11111000101101110010010011100000;
   assign mem[374175:374144] = 32'b11110110001110000010111011000000;
   assign mem[374207:374176] = 32'b00000010000101010011011011001000;
   assign mem[374239:374208] = 32'b00001000101111111000110011100000;
   assign mem[374271:374240] = 32'b11111100001010101101101110010000;
   assign mem[374303:374272] = 32'b00000001101001011101110001110110;
   assign mem[374335:374304] = 32'b00000101111101000001110010110000;
   assign mem[374367:374336] = 32'b11111001010000101110011001111000;
   assign mem[374399:374368] = 32'b00000111110110000100100000000000;
   assign mem[374431:374400] = 32'b11110110011010101100001101110000;
   assign mem[374463:374432] = 32'b11111111011010010001100011010100;
   assign mem[374495:374464] = 32'b11111101010011010100011000001000;
   assign mem[374527:374496] = 32'b00001000110000001010010100000000;
   assign mem[374559:374528] = 32'b11111100011011010100101110010000;
   assign mem[374591:374560] = 32'b00000001110011011001010011000100;
   assign mem[374623:374592] = 32'b00000001101001001010110010111100;
   assign mem[374655:374624] = 32'b11111010110111100000111110001000;
   assign mem[374687:374656] = 32'b00001011001010111100101000100000;
   assign mem[374719:374688] = 32'b11110010001110010110011001100000;
   assign mem[374751:374720] = 32'b11111011010001010010101000101000;
   assign mem[374783:374752] = 32'b11110111110111100111000000100000;
   assign mem[374815:374784] = 32'b00000010101101110000100010010000;
   assign mem[374847:374816] = 32'b00000100001000101010001010100000;
   assign mem[374879:374848] = 32'b11111110111010000100101001100000;
   assign mem[374911:374880] = 32'b11111111110000010000001110101000;
   assign mem[374943:374912] = 32'b00000001010011011101111010000100;
   assign mem[374975:374944] = 32'b11111000101101010111010100011000;
   assign mem[375007:374976] = 32'b00000011001111000111100100001100;
   assign mem[375039:375008] = 32'b11111101111101000101011111011000;
   assign mem[375071:375040] = 32'b00000010100011100100011000110000;
   assign mem[375103:375072] = 32'b11111110000110010000010100001010;
   assign mem[375135:375104] = 32'b00000000110100110000010001011010;
   assign mem[375167:375136] = 32'b11111101101010111110101111000100;
   assign mem[375199:375168] = 32'b00000010101110011010001101100100;
   assign mem[375231:375200] = 32'b11111011000011011100001001000000;
   assign mem[375263:375232] = 32'b11111100001100101110100110111100;
   assign mem[375295:375264] = 32'b00000011010001000100101000100000;
   assign mem[375327:375296] = 32'b11110111100010101000010110110000;
   assign mem[375359:375328] = 32'b00000001111110011111101110011010;
   assign mem[375391:375360] = 32'b00000011001000000010100110011000;
   assign mem[375423:375392] = 32'b00000011000000001100011010011100;
   assign mem[375455:375424] = 32'b00000001110101101000011111000000;
   assign mem[375487:375456] = 32'b11111111100100101100000010101010;
   assign mem[375519:375488] = 32'b00000010100010001111111011100000;
   assign mem[375551:375520] = 32'b00000010111010000000100000101000;
   assign mem[375583:375552] = 32'b00000001100010010011001000011110;
   assign mem[375615:375584] = 32'b11111101010001111001001000101100;
   assign mem[375647:375616] = 32'b00000000111110010100101001001000;
   assign mem[375679:375648] = 32'b11111101111111010001100111100000;
   assign mem[375711:375680] = 32'b00000110001100000000100101011000;
   assign mem[375743:375712] = 32'b11101111100101010011100010000000;
   assign mem[375775:375744] = 32'b00000101010010000100101000100000;
   assign mem[375807:375776] = 32'b00000100100011111100101000111000;
   assign mem[375839:375808] = 32'b00000001101010100000111011110000;
   assign mem[375871:375840] = 32'b11111110101000000101001100000000;
   assign mem[375903:375872] = 32'b00000011110011111100100111111000;
   assign mem[375935:375904] = 32'b11111111001111111000011010001100;
   assign mem[375967:375936] = 32'b00000000110101000000111001100010;
   assign mem[375999:375968] = 32'b00000010010101101000100010100100;
   assign mem[376031:376000] = 32'b11111010110000101001011011000000;
   assign mem[376063:376032] = 32'b00001000110111010001000100100000;
   assign mem[376095:376064] = 32'b00000000011101111010010110000101;
   assign mem[376127:376096] = 32'b00000001001100001011111000110010;
   assign mem[376159:376128] = 32'b11111101100100010001011010110100;
   assign mem[376191:376160] = 32'b00000000111100001001110011111010;
   assign mem[376223:376192] = 32'b11111111010000010111101101100111;
   assign mem[376255:376224] = 32'b11111001001001001101010000101000;
   assign mem[376287:376256] = 32'b11111111110101100000101000000001;
   assign mem[376319:376288] = 32'b00000000110100101001001100111010;
   assign mem[376351:376320] = 32'b00000000110100111000110111000000;
   assign mem[376383:376352] = 32'b00000011001010011001101101101100;
   assign mem[376415:376384] = 32'b11111000000000001011101000001000;
   assign mem[376447:376416] = 32'b00000010000001011110111011011000;
   assign mem[376479:376448] = 32'b11111111010011001100000001101000;
   assign mem[376511:376480] = 32'b00000010000011111000001101000100;
   assign mem[376543:376512] = 32'b00000001000101011101010111001100;
   assign mem[376575:376544] = 32'b11111110100110101001011011010110;
   assign mem[376607:376576] = 32'b00000001101111000011011111010010;
   assign mem[376639:376608] = 32'b00000000110110001000100110100111;
   assign mem[376671:376640] = 32'b11111011010111101110101011010000;
   assign mem[376703:376672] = 32'b00000010011011011110010000100000;
   assign mem[376735:376704] = 32'b00000000110000111010011101001100;
   assign mem[376767:376736] = 32'b00000000011000110100100000100100;
   assign mem[376799:376768] = 32'b00000001010100101101001010111110;
   assign mem[376831:376800] = 32'b00000010000010101111011101000100;
   assign mem[376863:376832] = 32'b11111101001100111101001100010000;
   assign mem[376895:376864] = 32'b00000001010000110001010011100110;
   assign mem[376927:376896] = 32'b00000001111010100000110100101110;
   assign mem[376959:376928] = 32'b00000010101100101111011101101100;
   assign mem[376991:376960] = 32'b11111101100111000101011011001100;
   assign mem[377023:376992] = 32'b00000001100110010101010000111110;
   assign mem[377055:377024] = 32'b11111100111110010001111110000100;
   assign mem[377087:377056] = 32'b11111101110010110001001111001100;
   assign mem[377119:377088] = 32'b11111110000100000010111011010110;
   assign mem[377151:377120] = 32'b11111010000111010010101011010000;
   assign mem[377183:377152] = 32'b11111111001110010111101100101011;
   assign mem[377215:377184] = 32'b11111110100001010010001101001000;
   assign mem[377247:377216] = 32'b00000010100000111001011000111000;
   assign mem[377279:377248] = 32'b11111111001000110111111011011010;
   assign mem[377311:377280] = 32'b00000101010110111010100101000000;
   assign mem[377343:377312] = 32'b00010010011011110110010100100000;
   assign mem[377375:377344] = 32'b00001110000001111011010011110000;
   assign mem[377407:377376] = 32'b11110011111001001101001100110000;
   assign mem[377439:377408] = 32'b11110111001000011001010001000000;
   assign mem[377471:377440] = 32'b00000010101010011110001001000100;
   assign mem[377503:377472] = 32'b11110001110111010011000001110000;
   assign mem[377535:377504] = 32'b00001001101110010001111010010000;
   assign mem[377567:377536] = 32'b11101110100001010011010101100000;
   assign mem[377599:377568] = 32'b00000010000110010010100010011000;
   assign mem[377631:377600] = 32'b11111011100001001001100101001000;
   assign mem[377663:377632] = 32'b11111101011111110010000100100000;
   assign mem[377695:377664] = 32'b00000001000001110001111100101100;
   assign mem[377727:377696] = 32'b11111111111100100001111110111101;
   assign mem[377759:377728] = 32'b00000101001111000111110110100000;
   assign mem[377791:377760] = 32'b11111011111111111100101011001000;
   assign mem[377823:377792] = 32'b00000101111111101111101101010000;
   assign mem[377855:377824] = 32'b00000001101110010000101111110000;
   assign mem[377887:377856] = 32'b00000000011011111010100010010000;
   assign mem[377919:377888] = 32'b11110100010100011110100100010000;
   assign mem[377951:377920] = 32'b00001001010110111110100110010000;
   assign mem[377983:377952] = 32'b11110011100110000010011111000000;
   assign mem[378015:377984] = 32'b00000110110001000110011101010000;
   assign mem[378047:378016] = 32'b11111011100011111011110001001000;
   assign mem[378079:378048] = 32'b11110111110010001100110110000000;
   assign mem[378111:378080] = 32'b00000001001010110110010110100100;
   assign mem[378143:378112] = 32'b00000100000110110101011100111000;
   assign mem[378175:378144] = 32'b11110011111101110001100000110000;
   assign mem[378207:378176] = 32'b11101111001101010111100000000000;
   assign mem[378239:378208] = 32'b11111101111010101011101100100000;
   assign mem[378271:378240] = 32'b00000010011000010101101011001100;
   assign mem[378303:378272] = 32'b00000001101110001001111010011100;
   assign mem[378335:378304] = 32'b11111110010100001101010111010000;
   assign mem[378367:378336] = 32'b00000000000110010111010001110011;
   assign mem[378399:378368] = 32'b00000001000000111010100100010010;
   assign mem[378431:378400] = 32'b00000000110100100001011100010011;
   assign mem[378463:378432] = 32'b11111011110010010111001000110000;
   assign mem[378495:378464] = 32'b00000010010101101010010010010000;
   assign mem[378527:378496] = 32'b11111100001011100010011111000000;
   assign mem[378559:378528] = 32'b00000010110001011000100100101100;
   assign mem[378591:378560] = 32'b00000011100000100101001100001100;
   assign mem[378623:378592] = 32'b11111011110001000010111100010000;
   assign mem[378655:378624] = 32'b11111110000110110010110010010000;
   assign mem[378687:378656] = 32'b11111100101011111000011111111100;
   assign mem[378719:378688] = 32'b00000100001111000010101000111000;
   assign mem[378751:378720] = 32'b11111110000001000110110110011110;
   assign mem[378783:378752] = 32'b00000011011100001010011010011100;
   assign mem[378815:378784] = 32'b00000110011001100000011000100000;
   assign mem[378847:378816] = 32'b11111111101111110101101001000001;
   assign mem[378879:378848] = 32'b11110111111101100100010111010000;
   assign mem[378911:378880] = 32'b11111100100000001100011110111000;
   assign mem[378943:378912] = 32'b11111010011101001100001011000000;
   assign mem[378975:378944] = 32'b00000100110011111010010001000000;
   assign mem[379007:378976] = 32'b00000110111000010001011001101000;
   assign mem[379039:379008] = 32'b11111110011110101110010101100010;
   assign mem[379071:379040] = 32'b11111101101111111001000001110000;
   assign mem[379103:379072] = 32'b00000100010101010101000010100000;
   assign mem[379135:379104] = 32'b11111111110011010110001101110110;
   assign mem[379167:379136] = 32'b11111101011010101101010100011000;
   assign mem[379199:379168] = 32'b11111011100011110111110110010000;
   assign mem[379231:379200] = 32'b00001000111001000101101110100000;
   assign mem[379263:379232] = 32'b00000000100010011100010011110111;
   assign mem[379295:379264] = 32'b00001000110011110101100110100000;
   assign mem[379327:379296] = 32'b11110111011101011010100100010000;
   assign mem[379359:379328] = 32'b00000000001100101110111100000100;
   assign mem[379391:379360] = 32'b00000011010011111101100101110000;
   assign mem[379423:379392] = 32'b00000100011111001001011000100000;
   assign mem[379455:379424] = 32'b00000001011110100010000001100000;
   assign mem[379487:379456] = 32'b11111010110100111110001110100000;
   assign mem[379519:379488] = 32'b11111100011011101111001111001100;
   assign mem[379551:379520] = 32'b11111010110010111111111100101000;
   assign mem[379583:379552] = 32'b11111111000011011111010011100101;
   assign mem[379615:379584] = 32'b00000000000111011010110010011101;
   assign mem[379647:379616] = 32'b00000000000100111110011100010000;
   assign mem[379679:379648] = 32'b00000101001011010100000001111000;
   assign mem[379711:379680] = 32'b11111010000010110011010000111000;
   assign mem[379743:379712] = 32'b00000000111100011101011001110110;
   assign mem[379775:379744] = 32'b00000110010000110111001101111000;
   assign mem[379807:379776] = 32'b00000001011011101100001000000010;
   assign mem[379839:379808] = 32'b11111010111011100100011001110000;
   assign mem[379871:379840] = 32'b00000001000011100101001011100110;
   assign mem[379903:379872] = 32'b00000011100000111010101111110100;
   assign mem[379935:379904] = 32'b00000000011000110101110000011101;
   assign mem[379967:379936] = 32'b11111110010011100000110100100010;
   assign mem[379999:379968] = 32'b11111100100100110111100110001100;
   assign mem[380031:380000] = 32'b00000001110110000110101011111000;
   assign mem[380063:380032] = 32'b11111101110111101100101110011000;
   assign mem[380095:380064] = 32'b00000011001100000011001010101100;
   assign mem[380127:380096] = 32'b11110101110110011101111001110000;
   assign mem[380159:380128] = 32'b00000011101100101011111110110100;
   assign mem[380191:380160] = 32'b00000000001101110100000001011011;
   assign mem[380223:380192] = 32'b11110111010000111111011000010000;
   assign mem[380255:380224] = 32'b00000001110110101110001000010010;
   assign mem[380287:380256] = 32'b00001000111011000000100101010000;
   assign mem[380319:380288] = 32'b11110010011010000011010001000000;
   assign mem[380351:380320] = 32'b00000110000010111101101010001000;
   assign mem[380383:380352] = 32'b00000001011001001100110110000010;
   assign mem[380415:380384] = 32'b11111011110101100000110001111000;
   assign mem[380447:380416] = 32'b00001001111111011000111100110000;
   assign mem[380479:380448] = 32'b11100001000110101001110110100000;
   assign mem[380511:380480] = 32'b11111100010110111010110101001100;
   assign mem[380543:380512] = 32'b11111011000011101111101100110000;
   assign mem[380575:380544] = 32'b00000010011001100111001111010100;
   assign mem[380607:380576] = 32'b00000111110001100100111000000000;
   assign mem[380639:380608] = 32'b11111010001011100111110110001000;
   assign mem[380671:380640] = 32'b00000101010000111101001011100000;
   assign mem[380703:380672] = 32'b00001001001000001110001110010000;
   assign mem[380735:380704] = 32'b11111000010101101101010101100000;
   assign mem[380767:380736] = 32'b00000101000111100001011000111000;
   assign mem[380799:380768] = 32'b11101100011001111011111110000000;
   assign mem[380831:380800] = 32'b11110111110111010010011101000000;
   assign mem[380863:380832] = 32'b00000101000010110000010111110000;
   assign mem[380895:380864] = 32'b11111101001000100111110110010000;
   assign mem[380927:380896] = 32'b11111001110111110001101110101000;
   assign mem[380959:380928] = 32'b00001010011000111101011001010000;
   assign mem[380991:380960] = 32'b11111101110010111011011001000100;
   assign mem[381023:380992] = 32'b00000110110110101100011111011000;
   assign mem[381055:381024] = 32'b00000101000001100111010110101000;
   assign mem[381087:381056] = 32'b11111100010010000110010001110100;
   assign mem[381119:381088] = 32'b00000010101000010111010011111100;
   assign mem[381151:381120] = 32'b11111011010011000010011101010000;
   assign mem[381183:381152] = 32'b11110101110100010100000111010000;
   assign mem[381215:381184] = 32'b00000011000111111010111000010100;
   assign mem[381247:381216] = 32'b00000000000000011110011110010000;
   assign mem[381279:381248] = 32'b11110011100000111110101001000000;
   assign mem[381311:381280] = 32'b11111110111100001000011100010000;
   assign mem[381343:381312] = 32'b11111000101011010111101110001000;
   assign mem[381375:381344] = 32'b00000110101100101011100011101000;
   assign mem[381407:381376] = 32'b00000011110110001010110000101000;
   assign mem[381439:381408] = 32'b00000100100011111111001110011000;
   assign mem[381471:381440] = 32'b11111000111010100110000010010000;
   assign mem[381503:381472] = 32'b11111100010011111010110011101000;
   assign mem[381535:381504] = 32'b00000000100010110000000110110100;
   assign mem[381567:381536] = 32'b11111101110110000011010111010000;
   assign mem[381599:381568] = 32'b00000100010011100110101010010000;
   assign mem[381631:381600] = 32'b00000100011110001111101110110000;
   assign mem[381663:381632] = 32'b00000010100110100110000010010000;
   assign mem[381695:381664] = 32'b11111101110000011101000110010000;
   assign mem[381727:381696] = 32'b00000010101100011100011111110100;
   assign mem[381759:381728] = 32'b00000011110110000010111001100000;
   assign mem[381791:381760] = 32'b00000001110100111100100111101100;
   assign mem[381823:381792] = 32'b00001001011100101110000111010000;
   assign mem[381855:381824] = 32'b11111110000000110110001101111100;
   assign mem[381887:381856] = 32'b11111000101110111110011010111000;
   assign mem[381919:381888] = 32'b00000111010001110110111100010000;
   assign mem[381951:381920] = 32'b11110100101101100011110101010000;
   assign mem[381983:381952] = 32'b11111111001010101101100100001010;
   assign mem[382015:381984] = 32'b00000011011100001101110111000100;
   assign mem[382047:382016] = 32'b11111111010000010100010010100001;
   assign mem[382079:382048] = 32'b00001000110101100101110001010000;
   assign mem[382111:382080] = 32'b11111111101110011011010000000001;
   assign mem[382143:382112] = 32'b00001011101010101110101101110000;
   assign mem[382175:382144] = 32'b11111111001110000010110111111001;
   assign mem[382207:382176] = 32'b00000010111110101011100010110000;
   assign mem[382239:382208] = 32'b11111001001000101011001011010000;
   assign mem[382271:382240] = 32'b00000010011010001110110101010000;
   assign mem[382303:382272] = 32'b00000000000000100001010011011100;
   assign mem[382335:382304] = 32'b11111001100110111110110011001000;
   assign mem[382367:382336] = 32'b00000001100000001100101101100110;
   assign mem[382399:382368] = 32'b11110110100100111011110111100000;
   assign mem[382431:382400] = 32'b11111001000000110011010110101000;
   assign mem[382463:382432] = 32'b11111111101111010011100000110111;
   assign mem[382495:382464] = 32'b11111100101001000100011101101100;
   assign mem[382527:382496] = 32'b00000100000100100010101110110000;
   assign mem[382559:382528] = 32'b11111001111000110011011110111000;
   assign mem[382591:382560] = 32'b00000011110010100111000001001100;
   assign mem[382623:382592] = 32'b00000011111100001111111110010000;
   assign mem[382655:382624] = 32'b11111011000110001110111100110000;
   assign mem[382687:382656] = 32'b00000010101111110100110101000000;
   assign mem[382719:382688] = 32'b00000000011110010011111101110111;
   assign mem[382751:382720] = 32'b11111011100001010011010010010000;
   assign mem[382783:382752] = 32'b00001010100001100010110100100000;
   assign mem[382815:382784] = 32'b11111100010100001110010010001100;
   assign mem[382847:382816] = 32'b11111101100110010111000011110100;
   assign mem[382879:382848] = 32'b00000111100010111111111101101000;
   assign mem[382911:382880] = 32'b11111110111001011110011101011110;
   assign mem[382943:382912] = 32'b00000110110001000010010100011000;
   assign mem[382975:382944] = 32'b00000110000110001101101100011000;
   assign mem[383007:382976] = 32'b11111010011000110000000000011000;
   assign mem[383039:383008] = 32'b11111000001111110111001101010000;
   assign mem[383071:383040] = 32'b11110001110100010100110011100000;
   assign mem[383103:383072] = 32'b11110111100001010100011100110000;
   assign mem[383135:383104] = 32'b00001001011110000111000000000000;
   assign mem[383167:383136] = 32'b00000101010011010001110001101000;
   assign mem[383199:383168] = 32'b00000100100011101101101011001000;
   assign mem[383231:383200] = 32'b00001000010010011010001101000000;
   assign mem[383263:383232] = 32'b00000101010101000010001111110000;
   assign mem[383295:383264] = 32'b11110010101010010111011100110000;
   assign mem[383327:383296] = 32'b00000001010100011111100011011000;
   assign mem[383359:383328] = 32'b11111000100101001001100110110000;
   assign mem[383391:383360] = 32'b00000000101100111011001111111001;
   assign mem[383423:383392] = 32'b11110101101100111011000111000000;
   assign mem[383455:383424] = 32'b00000000001001111111001111110111;
   assign mem[383487:383456] = 32'b11111101100111100010001000100100;
   assign mem[383519:383488] = 32'b00000001010100101111101011101000;
   assign mem[383551:383520] = 32'b11111111000111000111101000010111;
   assign mem[383583:383552] = 32'b11111100011001010110110111110100;
   assign mem[383615:383584] = 32'b00000010010111011110101000010000;
   assign mem[383647:383616] = 32'b11111100000101111011000100000100;
   assign mem[383679:383648] = 32'b00000101101100010101101110001000;
   assign mem[383711:383680] = 32'b11111110011000110110111001101110;
   assign mem[383743:383712] = 32'b11111111111101001101110101011010;
   assign mem[383775:383744] = 32'b11111100101100100000100101010100;
   assign mem[383807:383776] = 32'b11111011101011101011111111100000;
   assign mem[383839:383808] = 32'b00000010010101011110110010111000;
   assign mem[383871:383840] = 32'b11111101100110110000100101010100;
   assign mem[383903:383872] = 32'b11111011101100100100111100100000;
   assign mem[383935:383904] = 32'b00000010100110101000101010111000;
   assign mem[383967:383936] = 32'b00000000101010100010110111100011;
   assign mem[383999:383968] = 32'b11111101001000100010010000100000;
   assign mem[384031:384000] = 32'b11111011001010100101010100010000;
   assign mem[384063:384032] = 32'b00000010110101011010111111001000;
   assign mem[384095:384064] = 32'b00000000001010111111010110100011;
   assign mem[384127:384096] = 32'b11111100110001101101110010000000;
   assign mem[384159:384128] = 32'b00000100111010001000001111110000;
   assign mem[384191:384160] = 32'b11111010101110101010000011011000;
   assign mem[384223:384192] = 32'b11111111100010010010100000110001;
   assign mem[384255:384224] = 32'b00000011010010000000010110011100;
   assign mem[384287:384256] = 32'b11111101000010100011011011001100;
   assign mem[384319:384288] = 32'b11111111000000111111000101001001;
   assign mem[384351:384320] = 32'b00000001110001010000011011011010;
   assign mem[384383:384352] = 32'b11110111111001111101011001010000;
   assign mem[384415:384384] = 32'b00001000010100010001111001110000;
   assign mem[384447:384416] = 32'b11111111100110110101110100011010;
   assign mem[384479:384448] = 32'b00000011001000100011110111110000;
   assign mem[384511:384480] = 32'b11111100010001001011010100010000;
   assign mem[384543:384512] = 32'b11111100011110101111011010100100;
   assign mem[384575:384544] = 32'b00001001111000011110010010010000;
   assign mem[384607:384576] = 32'b11110111010110111011010010100000;
   assign mem[384639:384608] = 32'b00000001111101000100101101000000;
   assign mem[384671:384640] = 32'b11111111110110100011101001100000;
   assign mem[384703:384672] = 32'b11110011100101110000111101010000;
   assign mem[384735:384704] = 32'b00000001111100011010010011010000;
   assign mem[384767:384736] = 32'b00000011001011010011101100001100;
   assign mem[384799:384768] = 32'b11111010111010010110010010011000;
   assign mem[384831:384800] = 32'b00000010001010000010101100111100;
   assign mem[384863:384832] = 32'b00000010001110100001111110001000;
   assign mem[384895:384864] = 32'b11110111011101110101111011110000;
   assign mem[384927:384896] = 32'b00000011001000110100101110001000;
   assign mem[384959:384928] = 32'b11111111101111101110010110110111;
   assign mem[384991:384960] = 32'b00000110011011011100010111010000;
   assign mem[385023:384992] = 32'b00000100101101010000001100110000;
   assign mem[385055:385024] = 32'b11110001101010010110011011000000;
   assign mem[385087:385056] = 32'b11111011111101110100110011001000;
   assign mem[385119:385088] = 32'b00000001101000100000010010111110;
   assign mem[385151:385120] = 32'b00000011011001110001110101111000;
   assign mem[385183:385152] = 32'b11111111111110011100111001111110;
   assign mem[385215:385184] = 32'b00001010110000111001011000100000;
   assign mem[385247:385216] = 32'b11110100101110000101101101110000;
   assign mem[385279:385248] = 32'b00000010011100110001000011111100;
   assign mem[385311:385280] = 32'b00000011101000000000011100101000;
   assign mem[385343:385312] = 32'b11111010000100111111001100001000;
   assign mem[385375:385344] = 32'b00000011110000010100001000001100;
   assign mem[385407:385376] = 32'b11111111001011010101000100100110;
   assign mem[385439:385408] = 32'b00000010111001000111001010101000;
   assign mem[385471:385440] = 32'b11111101110000000011111011110000;
   assign mem[385503:385472] = 32'b00000101110100010110011101101000;
   assign mem[385535:385504] = 32'b11111110101000000101110011011100;
   assign mem[385567:385536] = 32'b00000001010111001010011000000100;
   assign mem[385599:385568] = 32'b11111001000110011010110010111000;
   assign mem[385631:385600] = 32'b11111110111011010100110100010000;
   assign mem[385663:385632] = 32'b11111011010100111011110111111000;
   assign mem[385695:385664] = 32'b00000001110010101011110000010010;
   assign mem[385727:385696] = 32'b00000101000011111100011011111000;
   assign mem[385759:385728] = 32'b00000000110111100010001111000111;
   assign mem[385791:385760] = 32'b00000010100000000111001010001000;
   assign mem[385823:385792] = 32'b00000001011001101000111111111100;
   assign mem[385855:385824] = 32'b00000011001101111101101111010000;
   assign mem[385887:385856] = 32'b00000001100110101100110010111000;
   assign mem[385919:385888] = 32'b11110011001100011100100111000000;
   assign mem[385951:385920] = 32'b00000101010100000001101101010000;
   assign mem[385983:385952] = 32'b11110110111011011000010101010000;
   assign mem[386015:385984] = 32'b11111101100111101110110001110100;
   assign mem[386047:386016] = 32'b00000001011110001100111111100010;
   assign mem[386079:386048] = 32'b00000010001000100110101001000100;
   assign mem[386111:386080] = 32'b11111111010101010001010101110011;
   assign mem[386143:386112] = 32'b00000011000101100010000001000100;
   assign mem[386175:386144] = 32'b00000100110001101101100111000000;
   assign mem[386207:386176] = 32'b11111111011101011100001000101011;
   assign mem[386239:386208] = 32'b00000010100000010101011011111100;
   assign mem[386271:386240] = 32'b00000101111110110010110110110000;
   assign mem[386303:386272] = 32'b00000100101010111010111101000000;
   assign mem[386335:386304] = 32'b00000010011000111001010110101000;
   assign mem[386367:386336] = 32'b11111110001011100110100101000100;
   assign mem[386399:386368] = 32'b11111011001000100001111010111000;
   assign mem[386431:386400] = 32'b00000000001001010000100100000011;
   assign mem[386463:386432] = 32'b11111110000111101011010010101100;
   assign mem[386495:386464] = 32'b00000001111001100010001110110110;
   assign mem[386527:386496] = 32'b11111011100001001100000010010000;
   assign mem[386559:386528] = 32'b00000000000110000110101100000010;
   assign mem[386591:386560] = 32'b00000001010000001110110111101110;
   assign mem[386623:386592] = 32'b11111111000001100111111100011111;
   assign mem[386655:386624] = 32'b11111011101001111001100111101000;
   assign mem[386687:386656] = 32'b00000100011111001011010111000000;
   assign mem[386719:386688] = 32'b11111011110010010010001100110000;
   assign mem[386751:386720] = 32'b00000001000011010010110011010100;
   assign mem[386783:386752] = 32'b00001001110100001111101111010000;
   assign mem[386815:386784] = 32'b11111100100000001000110100101100;
   assign mem[386847:386816] = 32'b11111101111111111010010010110000;
   assign mem[386879:386848] = 32'b00000101100011111100100001010000;
   assign mem[386911:386880] = 32'b11111000011000011000100101011000;
   assign mem[386943:386912] = 32'b00000011111111100111010111100000;
   assign mem[386975:386944] = 32'b11111101001101001011110111011100;
   assign mem[387007:386976] = 32'b00000110011100011101011100101000;
   assign mem[387039:387008] = 32'b11111110100010000010100110000110;
   assign mem[387071:387040] = 32'b00000110000011101101100100100000;
   assign mem[387103:387072] = 32'b11111111111101110011000001100100;
   assign mem[387135:387104] = 32'b11111100101001110100100011100000;
   assign mem[387167:387136] = 32'b00000011010110110110100000111100;
   assign mem[387199:387168] = 32'b11111101010011001011101101000000;
   assign mem[387231:387200] = 32'b00001001100000010100000010100000;
   assign mem[387263:387232] = 32'b00000001000000111101110011000100;
   assign mem[387295:387264] = 32'b11111111000000111101100011100001;
   assign mem[387327:387296] = 32'b11111010110100100000111101101000;
   assign mem[387359:387328] = 32'b11101101100000001001110010100000;
   assign mem[387391:387360] = 32'b00000100111000011110100111001000;
   assign mem[387423:387392] = 32'b00000011011100011011110000101000;
   assign mem[387455:387424] = 32'b11111110110010101011011011000000;
   assign mem[387487:387456] = 32'b11111000101100001000001011001000;
   assign mem[387519:387488] = 32'b11110100111100101101010001100000;
   assign mem[387551:387520] = 32'b11111111011001001111010000000010;
   assign mem[387583:387552] = 32'b11111111111101000000010111110010;
   assign mem[387615:387584] = 32'b00000001111010011010110011010000;
   assign mem[387647:387616] = 32'b00000000000101110110100001101100;
   assign mem[387679:387648] = 32'b11111100000000111010101011010000;
   assign mem[387711:387680] = 32'b00000011100000100010101011110100;
   assign mem[387743:387712] = 32'b00000011000010010010100000100000;
   assign mem[387775:387744] = 32'b11111010001111100000100110101000;
   assign mem[387807:387776] = 32'b00000001110000111000101000110100;
   assign mem[387839:387808] = 32'b11111000111011000110101001110000;
   assign mem[387871:387840] = 32'b00000001000010111100111001011100;
   assign mem[387903:387872] = 32'b11110100000110001111000110100000;
   assign mem[387935:387904] = 32'b00001010111001010100100011010000;
   assign mem[387967:387936] = 32'b00000010011010010010111100011000;
   assign mem[387999:387968] = 32'b11110101110110110110111110000000;
   assign mem[388031:388000] = 32'b11111111000010110110111100101011;
   assign mem[388063:388032] = 32'b11111100101100110011011000010000;
   assign mem[388095:388064] = 32'b00001001001000110010001110110000;
   assign mem[388127:388096] = 32'b00000010000010100110010100001000;
   assign mem[388159:388128] = 32'b00000011011111011001110111100000;
   assign mem[388191:388160] = 32'b00000100010110110100100001001000;
   assign mem[388223:388192] = 32'b11111000010001111111011111010000;
   assign mem[388255:388224] = 32'b00000011100111100110101001011000;
   assign mem[388287:388256] = 32'b11111010010011111010011000110000;
   assign mem[388319:388288] = 32'b11111100100101001010000000101000;
   assign mem[388351:388320] = 32'b11111111100001011001100111010100;
   assign mem[388383:388352] = 32'b00000000101100110001110001100011;
   assign mem[388415:388384] = 32'b00000111011110010110011101111000;
   assign mem[388447:388416] = 32'b11111000101011011110001101011000;
   assign mem[388479:388448] = 32'b11111101000111111100110001000000;
   assign mem[388511:388480] = 32'b00000010110110111001101011010000;
   assign mem[388543:388512] = 32'b00001000111110111001011001000000;
   assign mem[388575:388544] = 32'b00000001100111010010001011101000;
   assign mem[388607:388576] = 32'b11110100011110111110111001000000;
   assign mem[388639:388608] = 32'b11111110101110100110001110101110;
   assign mem[388671:388640] = 32'b11111010000001010100001001000000;
   assign mem[388703:388672] = 32'b11110111100011101000110011000000;
   assign mem[388735:388704] = 32'b00001010011101001011011101100000;
   assign mem[388767:388736] = 32'b11110001111010100000111000110000;
   assign mem[388799:388768] = 32'b00000001011000000101001101110010;
   assign mem[388831:388800] = 32'b00000010010001101111011011001100;
   assign mem[388863:388832] = 32'b00000010000001101010110110101000;
   assign mem[388895:388864] = 32'b00000010001011010111111100111000;
   assign mem[388927:388896] = 32'b00000001011001011001100111111100;
   assign mem[388959:388928] = 32'b11111101110110110001001100110100;
   assign mem[388991:388960] = 32'b11111100101010011110001100010000;
   assign mem[389023:388992] = 32'b11111101111101010101000111011100;
   assign mem[389055:389024] = 32'b00000011001011011010110100010000;
   assign mem[389087:389056] = 32'b11111001000110110100110010100000;
   assign mem[389119:389088] = 32'b11111111100000100011101111001001;
   assign mem[389151:389120] = 32'b00000001111111101011110110011000;
   assign mem[389183:389152] = 32'b00000010010100011100011101101100;
   assign mem[389215:389184] = 32'b00000101010110110011111001100000;
   assign mem[389247:389216] = 32'b11111101001011110111100000011100;
   assign mem[389279:389248] = 32'b11110100000001100110010010010000;
   assign mem[389311:389280] = 32'b11110110101000010101111000100000;
   assign mem[389343:389312] = 32'b00000001100011101110000010110010;
   assign mem[389375:389344] = 32'b00000101000000001100011001010000;
   assign mem[389407:389376] = 32'b11111100000110110001000111100000;
   assign mem[389439:389408] = 32'b11111101101000000101011101111100;
   assign mem[389471:389440] = 32'b11111001111000100100000000011000;
   assign mem[389503:389472] = 32'b11111101011000011010011010010000;
   assign mem[389535:389504] = 32'b11111100110011000010011100000000;
   assign mem[389567:389536] = 32'b00000100000111111010110010000000;
   assign mem[389599:389568] = 32'b11110111111011101010000000010000;
   assign mem[389631:389600] = 32'b00000010110011011000001100110100;
   assign mem[389663:389632] = 32'b00001000111110100011100101000000;
   assign mem[389695:389664] = 32'b11111001001100001101010111000000;
   assign mem[389727:389696] = 32'b00000100000000001101000011000000;
   assign mem[389759:389728] = 32'b11111011001101101101111001001000;
   assign mem[389791:389760] = 32'b11111011000010110101100110111000;
   assign mem[389823:389792] = 32'b11111011100001110000000111001000;
   assign mem[389855:389824] = 32'b00000011110000100110111111100100;
   assign mem[389887:389856] = 32'b00000000111000111001011111001000;
   assign mem[389919:389888] = 32'b11111101010111111000101000100000;
   assign mem[389951:389920] = 32'b00000100001111111100010111010000;
   assign mem[389983:389952] = 32'b00000010101011100010010010001100;
   assign mem[390015:389984] = 32'b11111000110010001000011100101000;
   assign mem[390047:390016] = 32'b00000101001000000001101100110000;
   assign mem[390079:390048] = 32'b00000000000110111011000101001101;
   assign mem[390111:390080] = 32'b00000000111000100110100001010011;
   assign mem[390143:390112] = 32'b11111010101000011100010001001000;
   assign mem[390175:390144] = 32'b00001101010010101010000101000000;
   assign mem[390207:390176] = 32'b11110110001111001111010000000000;
   assign mem[390239:390208] = 32'b00000100101110001110010010110000;
   assign mem[390271:390240] = 32'b11111010100000011011010011000000;
   assign mem[390303:390272] = 32'b11111011101001011110011001000000;
   assign mem[390335:390304] = 32'b00000110110001010011101101000000;
   assign mem[390367:390336] = 32'b11111110111110111100001111110100;
   assign mem[390399:390368] = 32'b11101100111011000000101110000000;
   assign mem[390431:390400] = 32'b00001011110101011101001010010000;
   assign mem[390463:390432] = 32'b00000000001001110111111001011111;
   assign mem[390495:390464] = 32'b00001010111111000110101011100000;
   assign mem[390527:390496] = 32'b11101011000000100000011000000000;
   assign mem[390559:390528] = 32'b00000100000010111100011100000000;
   assign mem[390591:390560] = 32'b11110111110000100110101100100000;
   assign mem[390623:390592] = 32'b11111011000000011100110011100000;
   assign mem[390655:390624] = 32'b11111111110101001011111110101000;
   assign mem[390687:390656] = 32'b00000010110001000011110101100000;
   assign mem[390719:390688] = 32'b11111010110011110001100110101000;
   assign mem[390751:390720] = 32'b00000011001010011011001011110000;
   assign mem[390783:390752] = 32'b11111010100101101101001011001000;
   assign mem[390815:390784] = 32'b00000010111011001010011000110100;
   assign mem[390847:390816] = 32'b00000000001001001101001100100011;
   assign mem[390879:390848] = 32'b00000001011011101000011001010000;
   assign mem[390911:390880] = 32'b11111101000000100011010001010000;
   assign mem[390943:390912] = 32'b00000000001101011011101011111100;
   assign mem[390975:390944] = 32'b00000101110000100100010011111000;
   assign mem[391007:390976] = 32'b11110010000010101101100100010000;
   assign mem[391039:391008] = 32'b11111110111111000110000011001100;
   assign mem[391071:391040] = 32'b00000100000000000110000001110000;
   assign mem[391103:391072] = 32'b11111101100000000000011101100000;
   assign mem[391135:391104] = 32'b11111111010101001110010000110001;
   assign mem[391167:391136] = 32'b00000010000001111011110010000000;
   assign mem[391199:391168] = 32'b00000001000001110110000010010100;
   assign mem[391231:391200] = 32'b11111101000111100001101000111100;
   assign mem[391263:391232] = 32'b11111111110011100010000001101110;
   assign mem[391295:391264] = 32'b00000001110011001100011101001010;
   assign mem[391327:391296] = 32'b00000001110001100100110011110110;
   assign mem[391359:391328] = 32'b00000001111011011100010011110110;
   assign mem[391391:391360] = 32'b00000101110001111110010111001000;
   assign mem[391423:391392] = 32'b11111110110100010100110101011000;
   assign mem[391455:391424] = 32'b00000001110000000110001010000000;
   assign mem[391487:391456] = 32'b11111010100101111110111010111000;
   assign mem[391519:391488] = 32'b11111010000011101111000010110000;
   assign mem[391551:391520] = 32'b11110101100011011011000010000000;
   assign mem[391583:391552] = 32'b00000101101110110001000101110000;
   assign mem[391615:391584] = 32'b00000010000101110010111001110000;
   assign mem[391647:391616] = 32'b00000000001111110010000001101001;
   assign mem[391679:391648] = 32'b11111110110000111010111101110000;
   assign mem[391711:391680] = 32'b11110111100111001100100100100000;
   assign mem[391743:391712] = 32'b00000101001011111010110010000000;
   assign mem[391775:391744] = 32'b00000100010100011111000101001000;
   assign mem[391807:391776] = 32'b11110111111111101101001100110000;
   assign mem[391839:391808] = 32'b11111111101110000011000100010101;
   assign mem[391871:391840] = 32'b00000110000000101011010001011000;
   assign mem[391903:391872] = 32'b11111111101000101101111100110110;
   assign mem[391935:391904] = 32'b00000110000010110100001011101000;
   assign mem[391967:391936] = 32'b00000000010001001111001001011110;
   assign mem[391999:391968] = 32'b11110010101111001000010010000000;
   assign mem[392031:392000] = 32'b00000010111100001101011001010000;
   assign mem[392063:392032] = 32'b11111101111110110110110111100000;
   assign mem[392095:392064] = 32'b11110001010010010110111000000000;
   assign mem[392127:392096] = 32'b00000000111001100111001010010001;
   assign mem[392159:392128] = 32'b00000000010001110010111001101101;
   assign mem[392191:392160] = 32'b11110110111010110100001000100000;
   assign mem[392223:392192] = 32'b00001011010010000001101100010000;
   assign mem[392255:392224] = 32'b00000011000101001001011111001000;
   assign mem[392287:392256] = 32'b11111000000000001011001001101000;
   assign mem[392319:392288] = 32'b00000110110000110111000110010000;
   assign mem[392351:392320] = 32'b00000001010110111000000101011110;
   assign mem[392383:392352] = 32'b00000001111011110000011101110000;
   assign mem[392415:392384] = 32'b00000110001101101111100101011000;
   assign mem[392447:392416] = 32'b11110001011111011110011000100000;
   assign mem[392479:392448] = 32'b00001001001101001010010111110000;
   assign mem[392511:392480] = 32'b11110111100100100010100100010000;
   assign mem[392543:392512] = 32'b11110011101011010010001011110000;
   assign mem[392575:392544] = 32'b00000101001000110100111101000000;
   assign mem[392607:392576] = 32'b11110100010111001001010011110000;
   assign mem[392639:392608] = 32'b11110101110011111110100101010000;
   assign mem[392671:392640] = 32'b11111111010111111110001011111011;
   assign mem[392703:392672] = 32'b11110100000001000101111101100000;
   assign mem[392735:392704] = 32'b00000110011011000110110111001000;
   assign mem[392767:392736] = 32'b00000000111000010110000100010010;
   assign mem[392799:392768] = 32'b00000100100100010011001110011000;
   assign mem[392831:392800] = 32'b11111101000111111101011000010000;
   assign mem[392863:392832] = 32'b11111100011011001101111011111100;
   assign mem[392895:392864] = 32'b11111000111110111010001110010000;
   assign mem[392927:392896] = 32'b00000010010010111001110100000100;
   assign mem[392959:392928] = 32'b11111011011010111111001000101000;
   assign mem[392991:392960] = 32'b11101101111110000110100110100000;
   assign mem[393023:392992] = 32'b00000110011111000100010000000000;
   assign mem[393055:393024] = 32'b00001100111101000010110011000000;
   assign mem[393087:393056] = 32'b11111000001001000100011000111000;
   assign mem[393119:393088] = 32'b00001010100101000100110111100000;
   assign mem[393151:393120] = 32'b11111011100011010110010101100000;
   assign mem[393183:393152] = 32'b11111000011100111100101010010000;
   assign mem[393215:393184] = 32'b00001010010100010010000010110000;
   assign mem[393247:393216] = 32'b11110101000110010100111001100000;
   assign mem[393279:393248] = 32'b00000000001001111011011100101011;
   assign mem[393311:393280] = 32'b11100001100101011001110100100000;
   assign mem[393343:393312] = 32'b00000011100100000101100010111000;
   assign mem[393375:393344] = 32'b00000011010100011011010101101000;
   assign mem[393407:393376] = 32'b11111110001101011000101100011100;
   assign mem[393439:393408] = 32'b00000011110001000011011110000000;
   assign mem[393471:393440] = 32'b11111101000000111011111000010100;
   assign mem[393503:393472] = 32'b11111110110001011110110101111110;
   assign mem[393535:393504] = 32'b00000110110100110010000000110000;
   assign mem[393567:393536] = 32'b11111111000100101011000100111101;
   assign mem[393599:393568] = 32'b11110111010111001010011010110000;
   assign mem[393631:393600] = 32'b11110111101010101001101000110000;
   assign mem[393663:393632] = 32'b00000000101101000111010111101110;
   assign mem[393695:393664] = 32'b00000101011111110010000000110000;
   assign mem[393727:393696] = 32'b00000010100101101111100001000000;
   assign mem[393759:393728] = 32'b00000110011110010101110010100000;
   assign mem[393791:393760] = 32'b11111101000101111011110101011100;
   assign mem[393823:393792] = 32'b11111110000010011101000100111010;
   assign mem[393855:393824] = 32'b00000100110110110110111100111000;
   assign mem[393887:393856] = 32'b00000000111001010001010101000101;
   assign mem[393919:393888] = 32'b00000001111111011010111000000000;
   assign mem[393951:393920] = 32'b00000101001000010111010111000000;
   assign mem[393983:393952] = 32'b11110111100011100001101001000000;
   assign mem[394015:393984] = 32'b11110010110000001111101100000000;
   assign mem[394047:394016] = 32'b11111100111100001001110010001100;
   assign mem[394079:394048] = 32'b11111001100110011000110110110000;
   assign mem[394111:394080] = 32'b11111100100010110001100010100100;
   assign mem[394143:394112] = 32'b00000000111000001110100110010000;
   assign mem[394175:394144] = 32'b00000110001001000110100101100000;
   assign mem[394207:394176] = 32'b00000000001010000101100110100111;
   assign mem[394239:394208] = 32'b11111001110110000000101010011000;
   assign mem[394271:394240] = 32'b00000100001011110101000111100000;
   assign mem[394303:394272] = 32'b11111011000010011111101001110000;
   assign mem[394335:394304] = 32'b00000011101001110010010110011100;
   assign mem[394367:394336] = 32'b11110111010100010110011000010000;
   assign mem[394399:394368] = 32'b00000000111011001100011000111101;
   assign mem[394431:394400] = 32'b11101111010011111100110010000000;
   assign mem[394463:394432] = 32'b00001000001010100011001001100000;
   assign mem[394495:394464] = 32'b00000101101000110100101111001000;
   assign mem[394527:394496] = 32'b11111011100110011100001110000000;
   assign mem[394559:394528] = 32'b11110100001010001111010101010000;
   assign mem[394591:394560] = 32'b11111011111001000000111110101000;
   assign mem[394623:394592] = 32'b11111011000111111101001100101000;
   assign mem[394655:394624] = 32'b11111011000111101100111111101000;
   assign mem[394687:394656] = 32'b00001000001111110111011000010000;
   assign mem[394719:394688] = 32'b00001010100111010011000111010000;
   assign mem[394751:394720] = 32'b11111110000101111100000001100110;
   assign mem[394783:394752] = 32'b11111110010011110110100000000100;
   assign mem[394815:394784] = 32'b00000010110110110100110001000000;
   assign mem[394847:394816] = 32'b11111111101111011101010111000001;
   assign mem[394879:394848] = 32'b11111111010011101111011111001000;
   assign mem[394911:394880] = 32'b11110101100100010001110010100000;
   assign mem[394943:394912] = 32'b00000000000000100100101001000101;
   assign mem[394975:394944] = 32'b00000010000110111100111101101000;
   assign mem[395007:394976] = 32'b11111100110011011001110101010000;
   assign mem[395039:395008] = 32'b00000100011010110111001111110000;
   assign mem[395071:395040] = 32'b11111010111001110100110111001000;
   assign mem[395103:395072] = 32'b11111110100111011100101111101010;
   assign mem[395135:395104] = 32'b00000100100001101101111010100000;
   assign mem[395167:395136] = 32'b00000010110010100001111001010000;
   assign mem[395199:395168] = 32'b11111001011100110001110011100000;
   assign mem[395231:395200] = 32'b00001001011111110011001100010000;
   assign mem[395263:395232] = 32'b00000000110100101011011111011111;
   assign mem[395295:395264] = 32'b00000001000111101110010011111000;
   assign mem[395327:395296] = 32'b11111110111011000111000000110010;
   assign mem[395359:395328] = 32'b11111111010010100110010100010001;
   assign mem[395391:395360] = 32'b11111000101001001010101100111000;
   assign mem[395423:395392] = 32'b00000011011101111100101010111100;
   assign mem[395455:395424] = 32'b11111111011100010110111101011101;
   assign mem[395487:395456] = 32'b00000101101001000110111101111000;
   assign mem[395519:395488] = 32'b11110101000100001001100110110000;
   assign mem[395551:395520] = 32'b00000100011100010000101010010000;
   assign mem[395583:395552] = 32'b11111100110111111101111101001100;
   assign mem[395615:395584] = 32'b00000011000111000111001010011100;
   assign mem[395647:395616] = 32'b11111001100111100010001111110000;
   assign mem[395679:395648] = 32'b00000001011110001101100100011100;
   assign mem[395711:395680] = 32'b11111101101101001001011010111100;
   assign mem[395743:395712] = 32'b11110111010110011110000011100000;
   assign mem[395775:395744] = 32'b00000101101000111010111111011000;
   assign mem[395807:395776] = 32'b11111010001101000101110011110000;
   assign mem[395839:395808] = 32'b11111101111110101000111101111000;
   assign mem[395871:395840] = 32'b11111100100111011100000000101100;
   assign mem[395903:395872] = 32'b00000010111000111010011011110000;
   assign mem[395935:395904] = 32'b00000011011011111001110010001000;
   assign mem[395967:395936] = 32'b00000011000001101111101111110100;
   assign mem[395999:395968] = 32'b00000100010110101010111111011000;
   assign mem[396031:396000] = 32'b11111101101100000111100110011100;
   assign mem[396063:396032] = 32'b00000100110010110011110000110000;
   assign mem[396095:396064] = 32'b11111010110101111110110110011000;
   assign mem[396127:396096] = 32'b00000011101010011011010110111100;
   assign mem[396159:396128] = 32'b11101001000000110001100111100000;
   assign mem[396191:396160] = 32'b00000101000010010000000000001000;
   assign mem[396223:396192] = 32'b11111110111001100110010100100000;
   assign mem[396255:396224] = 32'b00000001010010000011011011000110;
   assign mem[396287:396256] = 32'b00000010000101101000010011111000;
   assign mem[396319:396288] = 32'b11110110001011001001010010000000;
   assign mem[396351:396320] = 32'b11111101101101111110110101111000;
   assign mem[396383:396352] = 32'b00000011110001100110100010011100;
   assign mem[396415:396384] = 32'b00000011100011101011110001110000;
   assign mem[396447:396416] = 32'b11111011111001010100010110011000;
   assign mem[396479:396448] = 32'b11111111010111010011100011111010;
   assign mem[396511:396480] = 32'b11111110100001000000001001110100;
   assign mem[396543:396512] = 32'b11111100110001101011110101101100;
   assign mem[396575:396544] = 32'b11111111110101000000110001111000;
   assign mem[396607:396576] = 32'b11111111010010000010011010111011;
   assign mem[396639:396608] = 32'b00000011111101101010101101000100;
   assign mem[396671:396640] = 32'b00000010100011100001010110010100;
   assign mem[396703:396672] = 32'b00000010000011100010011010110100;
   assign mem[396735:396704] = 32'b11110111110101101100101001000000;
   assign mem[396767:396736] = 32'b00000001000010111001101010111100;
   assign mem[396799:396768] = 32'b00000101001000110110111000010000;
   assign mem[396831:396800] = 32'b11111111101101000111001010111100;
   assign mem[396863:396832] = 32'b11111011111110000101010110011000;
   assign mem[396895:396864] = 32'b11111011010011100001100111111000;
   assign mem[396927:396896] = 32'b00000000111001110101010011011010;
   assign mem[396959:396928] = 32'b00000100010110110001110110001000;
   assign mem[396991:396960] = 32'b00000100100110001000010010010000;
   assign mem[397023:396992] = 32'b11111011101101101001100000111000;
   assign mem[397055:397024] = 32'b11110100101110100101101010010000;
   assign mem[397087:397056] = 32'b00000011111011100000001100100100;
   assign mem[397119:397088] = 32'b00000011000001110101100001011100;
   assign mem[397151:397120] = 32'b00000001001001000111101011001000;
   assign mem[397183:397152] = 32'b11111011111001100011110101001000;
   assign mem[397215:397184] = 32'b11111101101101101110111010111000;
   assign mem[397247:397216] = 32'b00000000111010000010101000111110;
   assign mem[397279:397248] = 32'b00000001101001101011000110000110;
   assign mem[397311:397280] = 32'b00000000010000010011110010110111;
   assign mem[397343:397312] = 32'b00000000010110010010101000000011;
   assign mem[397375:397344] = 32'b11111111001111011100110011110110;
   assign mem[397407:397376] = 32'b11111101011001110011001110001100;
   assign mem[397439:397408] = 32'b11111111110101110110110001011011;
   assign mem[397471:397440] = 32'b11111100101111000000010001011000;
   assign mem[397503:397472] = 32'b00000000110011011101001010011011;
   assign mem[397535:397504] = 32'b11111100101110111101101101100100;
   assign mem[397567:397536] = 32'b11111101001000110000011001011100;
   assign mem[397599:397568] = 32'b00000101010010000000101110000000;
   assign mem[397631:397600] = 32'b11111110000111100010011111011000;
   assign mem[397663:397632] = 32'b11111001000011000100101011011000;
   assign mem[397695:397664] = 32'b00000010011011000100101011110100;
   assign mem[397727:397696] = 32'b00000000101101001011100011100010;
   assign mem[397759:397728] = 32'b11111111110010010011001010010101;
   assign mem[397791:397760] = 32'b11111110101111010110100111011110;
   assign mem[397823:397792] = 32'b11111100111010001100001110001000;
   assign mem[397855:397824] = 32'b00000101101011100111111001011000;
   assign mem[397887:397856] = 32'b11111101101011100101000110011000;
   assign mem[397919:397888] = 32'b00000101010110111100110011010000;
   assign mem[397951:397920] = 32'b11110000101011110010001010100000;
   assign mem[397983:397952] = 32'b11110100010011111101000001100000;
   assign mem[398015:397984] = 32'b00000011010101100000000111001000;
   assign mem[398047:398016] = 32'b11111011111101000111100101001000;
   assign mem[398079:398048] = 32'b00000001011011101010101111100110;
   assign mem[398111:398080] = 32'b00000011100001001001010111010000;
   assign mem[398143:398112] = 32'b00000101011111011111100111101000;
   assign mem[398175:398144] = 32'b00001000001111001010100101100000;
   assign mem[398207:398176] = 32'b11111100101110110010110011001100;
   assign mem[398239:398208] = 32'b00000011001110111101110100111100;
   assign mem[398271:398240] = 32'b11110101101011110101001101010000;
   assign mem[398303:398272] = 32'b11111111110111011111000100011100;
   assign mem[398335:398304] = 32'b00000000011110111100000111101101;
   assign mem[398367:398336] = 32'b00000000111010010001010010111010;
   assign mem[398399:398368] = 32'b11110101100100110010100000000000;
   assign mem[398431:398400] = 32'b11111000101110001110010001100000;
   assign mem[398463:398432] = 32'b11111110000011000110101100000000;
   assign mem[398495:398464] = 32'b00000100110011011100010010001000;
   assign mem[398527:398496] = 32'b00000010001011110110010111000100;
   assign mem[398559:398528] = 32'b00000011011100100011100101110100;
   assign mem[398591:398560] = 32'b00000100101011110000000001001000;
   assign mem[398623:398592] = 32'b00000000110000000110110101101001;
   assign mem[398655:398624] = 32'b11111010100101001100101010110000;
   assign mem[398687:398656] = 32'b00000000100011110111101011110100;
   assign mem[398719:398688] = 32'b11110111001101110001100010010000;
   assign mem[398751:398720] = 32'b11111111000100001011001000110111;
   assign mem[398783:398752] = 32'b11111010011100101001101010011000;
   assign mem[398815:398784] = 32'b11111010101100010101011101011000;
   assign mem[398847:398816] = 32'b00000101010100011001000101001000;
   assign mem[398879:398848] = 32'b00000110101101010101101001000000;
   assign mem[398911:398880] = 32'b11111101100011101111101110010000;
   assign mem[398943:398912] = 32'b11111110101101100100000001110100;
   assign mem[398975:398944] = 32'b11111010110010001011001101110000;
   assign mem[399007:398976] = 32'b00000001101010101111100000110010;
   assign mem[399039:399008] = 32'b00000010000001000100001110010100;
   assign mem[399071:399040] = 32'b00000101111100000101010100100000;
   assign mem[399103:399072] = 32'b11110101010010101011001001110000;
   assign mem[399135:399104] = 32'b00001010101100101111011010110000;
   assign mem[399167:399136] = 32'b11110010111011000000101100110000;
   assign mem[399199:399168] = 32'b00000111010101001110000111010000;
   assign mem[399231:399200] = 32'b11110101010111000011111001110000;
   assign mem[399263:399232] = 32'b11111101100101011011011110000100;
   assign mem[399295:399264] = 32'b00000110010110100100000111111000;
   assign mem[399327:399296] = 32'b11111001111101110011101111010000;
   assign mem[399359:399328] = 32'b11110110100010011110110000000000;
   assign mem[399391:399360] = 32'b00000010111010111100100010110100;
   assign mem[399423:399392] = 32'b00000010001100111110011011010100;
   assign mem[399455:399424] = 32'b00000010111000101001110011011100;
   assign mem[399487:399456] = 32'b11111111101110001000110101101010;
   assign mem[399519:399488] = 32'b11111001000000100011000111011000;
   assign mem[399551:399520] = 32'b11111110000100110001001000101010;
   assign mem[399583:399552] = 32'b00000010101000101100000110000100;
   assign mem[399615:399584] = 32'b00000110001110111010111011001000;
   assign mem[399647:399616] = 32'b11111000000001101111011100011000;
   assign mem[399679:399648] = 32'b00000100100111111100100101101000;
   assign mem[399711:399680] = 32'b00001000110100100000001001110000;
   assign mem[399743:399712] = 32'b11101111001100111111001010100000;
   assign mem[399775:399744] = 32'b00001000101101010111110000110000;
   assign mem[399807:399776] = 32'b11111110100111100100100011010010;
   assign mem[399839:399808] = 32'b11111110011000110000011111101110;
   assign mem[399871:399840] = 32'b11111111001101111100000111110010;
   assign mem[399903:399872] = 32'b11111101100100100101100110110000;
   assign mem[399935:399904] = 32'b00001100100011010101010010010000;
   assign mem[399967:399936] = 32'b11110000001011011111110110100000;
   assign mem[399999:399968] = 32'b00000000100001110101011001000100;
   assign mem[400031:400000] = 32'b00000100011000110001010011000000;
   assign mem[400063:400032] = 32'b11111111001000011100000001101111;
   assign mem[400095:400064] = 32'b00000110101101010001001111100000;
   assign mem[400127:400096] = 32'b11111000111101110000100001011000;
   assign mem[400159:400128] = 32'b00000111101111010011101101111000;
   assign mem[400191:400160] = 32'b11111001011001010110110001000000;
   assign mem[400223:400192] = 32'b11111101110110001001100111100100;
   assign mem[400255:400224] = 32'b00000111010111110101100011011000;
   assign mem[400287:400256] = 32'b11111000011101100000101111001000;
   assign mem[400319:400288] = 32'b11111011011111000110101111001000;
   assign mem[400351:400320] = 32'b00000011001000010011110000111000;
   assign mem[400383:400352] = 32'b11111010011100010110001011101000;
   assign mem[400415:400384] = 32'b11111010101110110010100000001000;
   assign mem[400447:400416] = 32'b00000010111111110001011011000000;
   assign mem[400479:400448] = 32'b11111110011000001000110011011110;
   assign mem[400511:400480] = 32'b00000001011000001101000100001100;
   assign mem[400543:400512] = 32'b00000011000000010101111001011100;
   assign mem[400575:400544] = 32'b00000110001010011101010101101000;
   assign mem[400607:400576] = 32'b11111101100100011000000101110000;
   assign mem[400639:400608] = 32'b00000001000101011010101001111000;
   assign mem[400671:400640] = 32'b11110001000000000000011001010000;
   assign mem[400703:400672] = 32'b00000010010000001011111000001000;
   assign mem[400735:400704] = 32'b00000001111111010010011000010100;
   assign mem[400767:400736] = 32'b00000001100001010101011101000010;
   assign mem[400799:400768] = 32'b11111001101011111000110010110000;
   assign mem[400831:400800] = 32'b00000000001111101010001010010011;
   assign mem[400863:400832] = 32'b00000111000010100010000101011000;
   assign mem[400895:400864] = 32'b00000100011100111010111010110000;
   assign mem[400927:400896] = 32'b00001000001101110010110100000000;
   assign mem[400959:400928] = 32'b11101110100101100111100111000000;
   assign mem[400991:400960] = 32'b11110001010101111100010101100000;
   assign mem[401023:400992] = 32'b00000010011101000111111100100000;
   assign mem[401055:401024] = 32'b11111111001011100100010111100110;
   assign mem[401087:401056] = 32'b00000100010010110111010001110000;
   assign mem[401119:401088] = 32'b00000101011111100101110101010000;
   assign mem[401151:401120] = 32'b00000001100110110111010001010100;
   assign mem[401183:401152] = 32'b11111100101001111110000110100100;
   assign mem[401215:401184] = 32'b00001001000111000011101011000000;
   assign mem[401247:401216] = 32'b00000100101110111000100001101000;
   assign mem[401279:401248] = 32'b11111001110111010011001011100000;
   assign mem[401311:401280] = 32'b00000011010001100111111101010100;
   assign mem[401343:401312] = 32'b11111110001100001000000111011110;
   assign mem[401375:401344] = 32'b00000011001001101100011111101000;
   assign mem[401407:401376] = 32'b11111100000110010100101111101000;
   assign mem[401439:401408] = 32'b00000100100100100001011011100000;
   assign mem[401471:401440] = 32'b11111001011001000011111010101000;
   assign mem[401503:401472] = 32'b00000100011111111111000101111000;
   assign mem[401535:401504] = 32'b00000011101100111001111011001100;
   assign mem[401567:401536] = 32'b11110001011000111001110001010000;
   assign mem[401599:401568] = 32'b11111101010110100111001110011000;
   assign mem[401631:401600] = 32'b11111111111101110110010011011100;
   assign mem[401663:401632] = 32'b11111010001000110101010111011000;
   assign mem[401695:401664] = 32'b00001100010000010011111101000000;
   assign mem[401727:401696] = 32'b11101101010101011100111000100000;
   assign mem[401759:401728] = 32'b11111001111011110101110100100000;
   assign mem[401791:401760] = 32'b00000010100101001010100011011100;
   assign mem[401823:401792] = 32'b11101100111001000100011000000000;
   assign mem[401855:401824] = 32'b11111110100010010000100100111110;
   assign mem[401887:401856] = 32'b00000110001010101000111110101000;
   assign mem[401919:401888] = 32'b11111000100110010100101100101000;
   assign mem[401951:401920] = 32'b00000101010110100010111010101000;
   assign mem[401983:401952] = 32'b11110101000000111000110100100000;
   assign mem[402015:401984] = 32'b00001101000001100110101111010000;
   assign mem[402047:402016] = 32'b11111000110111111111011000110000;
   assign mem[402079:402048] = 32'b11111110010000100101010010110110;
   assign mem[402111:402080] = 32'b00000000011111101001111101010100;
   assign mem[402143:402112] = 32'b00000010110001000101001101011000;
   assign mem[402175:402144] = 32'b11111111101000111000111011111101;
   assign mem[402207:402176] = 32'b11111011101000011011100100110000;
   assign mem[402239:402208] = 32'b00000001101111011100011000011110;
   assign mem[402271:402240] = 32'b00001000101110101010110001010000;
   assign mem[402303:402272] = 32'b11110010110001001011101101110000;
   assign mem[402335:402304] = 32'b11111111000101001111100011000011;
   assign mem[402367:402336] = 32'b11110110110101001111111000100000;
   assign mem[402399:402368] = 32'b00000100110011001100001010111000;
   assign mem[402431:402400] = 32'b11101010000111010011010011100000;
   assign mem[402463:402432] = 32'b00000100000100110011111110111000;
   assign mem[402495:402464] = 32'b00001000101111000010001110010000;
   assign mem[402527:402496] = 32'b11111101100100000001101000000000;
   assign mem[402559:402528] = 32'b00000001001011010001010011111100;
   assign mem[402591:402560] = 32'b11111101000111000000010100001100;
   assign mem[402623:402592] = 32'b00000000011010011010001101111010;
   assign mem[402655:402624] = 32'b00010001000010011010010011000000;
   assign mem[402687:402656] = 32'b11101000000101011100101001100000;
   assign mem[402719:402688] = 32'b11111100011001100010111000010100;
   assign mem[402751:402720] = 32'b00000100110000110010011100101000;
   assign mem[402783:402752] = 32'b11110001110101101110101010100000;
   assign mem[402815:402784] = 32'b00000101011111000100011111011000;
   assign mem[402847:402816] = 32'b11111100100010011101100000110100;
   assign mem[402879:402848] = 32'b11111101000010100100010010111000;
   assign mem[402911:402880] = 32'b00000001100000110001110010110100;
   assign mem[402943:402912] = 32'b00000001010100101111011011111010;
   assign mem[402975:402944] = 32'b11111011100101101100111011000000;
   assign mem[403007:402976] = 32'b00000100001001001100111111101000;
   assign mem[403039:403008] = 32'b11111101000000001010101011010000;
   assign mem[403071:403040] = 32'b00000100101100101011011001000000;
   assign mem[403103:403072] = 32'b00000101110000110101100110100000;
   assign mem[403135:403104] = 32'b11111011110001101100110110100000;
   assign mem[403167:403136] = 32'b00000100010001101000000010110000;
   assign mem[403199:403168] = 32'b00000000001100110111100111110100;
   assign mem[403231:403200] = 32'b11111011111001010011011001010000;
   assign mem[403263:403232] = 32'b00000000010001111010010101000111;
   assign mem[403295:403264] = 32'b00000101111000010111101100110000;
   assign mem[403327:403296] = 32'b00000010100100010101001101011000;
   assign mem[403359:403328] = 32'b00000001001111011110000111010110;
   assign mem[403391:403360] = 32'b00000001010010100011010110000100;
   assign mem[403423:403392] = 32'b00000000000011010111011000110111;
   assign mem[403455:403424] = 32'b00000011110001101000011100110100;
   assign mem[403487:403456] = 32'b11101100101100000011001010100000;
   assign mem[403519:403488] = 32'b00000001100000100100110110011110;
   assign mem[403551:403520] = 32'b11111001110001110011000010100000;
   assign mem[403583:403552] = 32'b11111100101101100000001100111000;
   assign mem[403615:403584] = 32'b11111000100100110111011110010000;
   assign mem[403647:403616] = 32'b00000110111010110101100011101000;
   assign mem[403679:403648] = 32'b11110101000101000001111110110000;
   assign mem[403711:403680] = 32'b00001000010101111100001111110000;
   assign mem[403743:403712] = 32'b00000100011001011110001101000000;
   assign mem[403775:403744] = 32'b11111101110001100011000111000100;
   assign mem[403807:403776] = 32'b00000110000111100101101001100000;
   assign mem[403839:403808] = 32'b11111010011110111000111000101000;
   assign mem[403871:403840] = 32'b00000011111101110110111110000000;
   assign mem[403903:403872] = 32'b11111100100001100101111000011000;
   assign mem[403935:403904] = 32'b00000110000100110000100000111000;
   assign mem[403967:403936] = 32'b11111101100111010010001001011000;
   assign mem[403999:403968] = 32'b11111010011111000010111001000000;
   assign mem[404031:404000] = 32'b00000011011110000011111011010000;
   assign mem[404063:404032] = 32'b11111001001011111110100011010000;
   assign mem[404095:404064] = 32'b11111011111100010110111101100000;
   assign mem[404127:404096] = 32'b00000010001000101000011111011000;
   assign mem[404159:404128] = 32'b11110100110100101001101100010000;
   assign mem[404191:404160] = 32'b00000001001111010001011010010000;
   assign mem[404223:404192] = 32'b11111110010010110010000010110100;
   assign mem[404255:404224] = 32'b00000001011110110100001100001110;
   assign mem[404287:404256] = 32'b00000001011101001111111110001010;
   assign mem[404319:404288] = 32'b11111111100111001001000111101111;
   assign mem[404351:404320] = 32'b00000000000111110010111110000100;
   assign mem[404383:404352] = 32'b00000001011100111110010000001100;
   assign mem[404415:404384] = 32'b11111111011010111001011011000101;
   assign mem[404447:404416] = 32'b11111101011110100101010111111000;
   assign mem[404479:404448] = 32'b00000000001110110001110100101001;
   assign mem[404511:404480] = 32'b00000001100011011011110111000010;
   assign mem[404543:404512] = 32'b11111101011111111000000001101100;
   assign mem[404575:404544] = 32'b11111111000111110100101010011010;
   assign mem[404607:404576] = 32'b11111110000011111001000000101100;
   assign mem[404639:404608] = 32'b00000101100110101100111110001000;
   assign mem[404671:404640] = 32'b11111101110110010000100100101000;
   assign mem[404703:404672] = 32'b00000011001011101110111010010000;
   assign mem[404735:404704] = 32'b00000001111111000110010100111100;
   assign mem[404767:404736] = 32'b11110001111101101001011110010000;
   assign mem[404799:404768] = 32'b00000011000000101000111011100100;
   assign mem[404831:404800] = 32'b11111001000111011011001000101000;
   assign mem[404863:404832] = 32'b11111101110010110110000110110000;
   assign mem[404895:404864] = 32'b00001110011000011010110001000000;
   assign mem[404927:404896] = 32'b11111100101100100010111111100100;
   assign mem[404959:404928] = 32'b11111100110101010011000001110100;
   assign mem[404991:404960] = 32'b11111010100000110000011010101000;
   assign mem[405023:404992] = 32'b00000000000100100110010100001011;
   assign mem[405055:405024] = 32'b00001001001110101000100011000000;
   assign mem[405087:405056] = 32'b11110100100001110110000101000000;
   assign mem[405119:405088] = 32'b11111110010000101100010010111000;
   assign mem[405151:405120] = 32'b00000011010110101001000001111000;
   assign mem[405183:405152] = 32'b00000000000001100101111011111101;
   assign mem[405215:405184] = 32'b11111101011001000101011001011000;
   assign mem[405247:405216] = 32'b00000011001010101001010101000100;
   assign mem[405279:405248] = 32'b11111111111001101111110110111101;
   assign mem[405311:405280] = 32'b00000000001110111010001011110100;
   assign mem[405343:405312] = 32'b00000010101010100111010010111000;
   assign mem[405375:405344] = 32'b00000001100100001011100011001100;
   assign mem[405407:405376] = 32'b00000011000000111000010111001000;
   assign mem[405439:405408] = 32'b11111100110010100110000011100100;
   assign mem[405471:405440] = 32'b00000001011101010000000101010100;
   assign mem[405503:405472] = 32'b00001011111111011001010000110000;
   assign mem[405535:405504] = 32'b11101110110011111100111100000000;
   assign mem[405567:405536] = 32'b11111110110001101111111001100010;
   assign mem[405599:405568] = 32'b11110111100001101000110110000000;
   assign mem[405631:405600] = 32'b00000001010100010000010110001010;
   assign mem[405663:405632] = 32'b11111100010011111011100010010100;
   assign mem[405695:405664] = 32'b11111000010110000110011010101000;
   assign mem[405727:405696] = 32'b00001011010001010110111100110000;
   assign mem[405759:405728] = 32'b11111100110111000001100110001000;
   assign mem[405791:405760] = 32'b00001001101010001001101101110000;
   assign mem[405823:405792] = 32'b11111101001010000000001110000100;
   assign mem[405855:405824] = 32'b00000111110100000010101111101000;
   assign mem[405887:405856] = 32'b11110111001100110111010010000000;
   assign mem[405919:405888] = 32'b00000011111000011010101101101100;
   assign mem[405951:405920] = 32'b11111001111111011101011100111000;
   assign mem[405983:405952] = 32'b00000001101001000111101111110010;
   assign mem[406015:405984] = 32'b00000111011100000101000100011000;
   assign mem[406047:406016] = 32'b11111101111011011110011100001000;
   assign mem[406079:406048] = 32'b11101101110011100100110000000000;
   assign mem[406111:406080] = 32'b11111011000010110111011101101000;
   assign mem[406143:406112] = 32'b00000010101111100101000011100100;
   assign mem[406175:406144] = 32'b00000001110000000100101010000010;
   assign mem[406207:406176] = 32'b11111011101110010010000000011000;
   assign mem[406239:406208] = 32'b00000100010011111001101001000000;
   assign mem[406271:406240] = 32'b00000001111011011000110010001000;
   assign mem[406303:406272] = 32'b11111101110100010010101000010000;
   assign mem[406335:406304] = 32'b00000001011011100001010110001000;
   assign mem[406367:406336] = 32'b00000000100100001110101101100101;
   assign mem[406399:406368] = 32'b11101011111111111111100010000000;
   assign mem[406431:406400] = 32'b00000111110010011101011011110000;
   assign mem[406463:406432] = 32'b11111101000110001100100110110100;
   assign mem[406495:406464] = 32'b00000100010100111101101101100000;
   assign mem[406527:406496] = 32'b11111111000000111101010010011111;
   assign mem[406559:406528] = 32'b00000010000010010011101011010000;
   assign mem[406591:406560] = 32'b11111000100100101101001110100000;
   assign mem[406623:406592] = 32'b00000010111011110000100000110100;
   assign mem[406655:406624] = 32'b00000111001011000100110010111000;
   assign mem[406687:406656] = 32'b11111000101100100000001001110000;
   assign mem[406719:406688] = 32'b11111000001000101011010111011000;
   assign mem[406751:406720] = 32'b11111110101001111000101011111100;
   assign mem[406783:406752] = 32'b11101110110001001001001111000000;
   assign mem[406815:406784] = 32'b11111110101010111110100110000000;
   assign mem[406847:406816] = 32'b00000011100000001110100100001000;
   assign mem[406879:406848] = 32'b11110110111011011110101110110000;
   assign mem[406911:406880] = 32'b11111110000001101010011011010000;
   assign mem[406943:406912] = 32'b00000010010110000101111001010000;
   assign mem[406975:406944] = 32'b00000100011100010100101110111000;
   assign mem[407007:406976] = 32'b11111111111110100010110111100011;
   assign mem[407039:407008] = 32'b11111101001101101111101001010000;
   assign mem[407071:407040] = 32'b11111110110101100101000000010000;
   assign mem[407103:407072] = 32'b11111000100101001110001111100000;
   assign mem[407135:407104] = 32'b11111000001011110001100100101000;
   assign mem[407167:407136] = 32'b00000000110001000000101100011100;
   assign mem[407199:407168] = 32'b11111101100100100010011110101100;
   assign mem[407231:407200] = 32'b00000010010100110101101001011100;
   assign mem[407263:407232] = 32'b00000010000001111010101101111000;
   assign mem[407295:407264] = 32'b11111101110111000100011011010000;
   assign mem[407327:407296] = 32'b00000001100000100010011010100000;
   assign mem[407359:407328] = 32'b00000001001000110000010000000110;
   assign mem[407391:407360] = 32'b00000010000111000000111000101100;
   assign mem[407423:407392] = 32'b11111110001111110100110111010010;
   assign mem[407455:407424] = 32'b00000100110111001110010010010000;
   assign mem[407487:407456] = 32'b00000001111110000011010100011100;
   assign mem[407519:407488] = 32'b11111101010101110011010101100100;
   assign mem[407551:407520] = 32'b00000010111111100001010001011000;
   assign mem[407583:407552] = 32'b11111110011011111001000011011010;
   assign mem[407615:407584] = 32'b11111011010000010000010111010000;
   assign mem[407647:407616] = 32'b00000001010010111010011010011000;
   assign mem[407679:407648] = 32'b11110000001011100001010000110000;
   assign mem[407711:407680] = 32'b11110010110011000110000101010000;
   assign mem[407743:407712] = 32'b00000000000111111101101000110010;
   assign mem[407775:407744] = 32'b00000001111100000111101101111010;
   assign mem[407807:407776] = 32'b00001000110001100100001100110000;
   assign mem[407839:407808] = 32'b11101111010011010000010111100000;
   assign mem[407871:407840] = 32'b00000001001100010110100110111100;
   assign mem[407903:407872] = 32'b00000010000101001011010111001100;
   assign mem[407935:407904] = 32'b11111000000001110010001111011000;
   assign mem[407967:407936] = 32'b00000010110100000000111110011000;
   assign mem[407999:407968] = 32'b11111000101011010001100101000000;
   assign mem[408031:408000] = 32'b11111001001111110101000100001000;
   assign mem[408063:408032] = 32'b11111110000011010001101101001110;
   assign mem[408095:408064] = 32'b11111011101100011001011100001000;
   assign mem[408127:408096] = 32'b00000011101101101010101000101100;
   assign mem[408159:408128] = 32'b11111000101011100110010110011000;
   assign mem[408191:408160] = 32'b00000001110010010100100100100010;
   assign mem[408223:408192] = 32'b00000110000111111011110101111000;
   assign mem[408255:408224] = 32'b11110111011001110000110010100000;
   assign mem[408287:408256] = 32'b00000101111101100000000111111000;
   assign mem[408319:408288] = 32'b11111000010111101000001101011000;
   assign mem[408351:408320] = 32'b11110111010111000010111000110000;
   assign mem[408383:408352] = 32'b00000000100111111101100001101110;
   assign mem[408415:408384] = 32'b00010011110111110010110010100000;
   assign mem[408447:408416] = 32'b11110010110001000011111000010000;
   assign mem[408479:408448] = 32'b00000011001010000111110011001000;
   assign mem[408511:408480] = 32'b00000010110110101001100001110100;
   assign mem[408543:408512] = 32'b11111011110001111100010111001000;
   assign mem[408575:408544] = 32'b00001001011110010000010000010000;
   assign mem[408607:408576] = 32'b11110100110000010001110110010000;
   assign mem[408639:408608] = 32'b11111010011011110110110111101000;
   assign mem[408671:408640] = 32'b00000000101100011000001000111011;
   assign mem[408703:408672] = 32'b11111101100000110110010010010100;
   assign mem[408735:408704] = 32'b00010011010011010100001101000000;
   assign mem[408767:408736] = 32'b11111101110100100101001111100100;
   assign mem[408799:408768] = 32'b00001010000010000111110101000000;
   assign mem[408831:408800] = 32'b11111111011111101010111011000111;
   assign mem[408863:408832] = 32'b00000001000101000111101001001000;
   assign mem[408895:408864] = 32'b00001111111110100010111100010000;
   assign mem[408927:408896] = 32'b11110000010010000100100000010000;
   assign mem[408959:408928] = 32'b11111001010000100100101111110000;
   assign mem[408991:408960] = 32'b00000001101100101100000101000100;
   assign mem[409023:408992] = 32'b11111011111010010100110010010000;
   assign mem[409055:409024] = 32'b00000101101011100001011111010000;
   assign mem[409087:409056] = 32'b11110111111100010100000110000000;
   assign mem[409119:409088] = 32'b00000100001111100010001000010000;
   assign mem[409151:409120] = 32'b11111110100011110010110011000100;
   assign mem[409183:409152] = 32'b11111101000011000001110100010000;
   assign mem[409215:409184] = 32'b00000000101011001011010001011010;
   assign mem[409247:409216] = 32'b11110010000000101001001110110000;
   assign mem[409279:409248] = 32'b00000110011011111101111101010000;
   assign mem[409311:409280] = 32'b00001000111011000100011101100000;
   assign mem[409343:409312] = 32'b11110001010010000011011001110000;
   assign mem[409375:409344] = 32'b11110111001011110111000101010000;
   assign mem[409407:409376] = 32'b11111101111100010100000111111000;
   assign mem[409439:409408] = 32'b11111111101110001001010110110011;
   assign mem[409471:409440] = 32'b11111110100000101001011100100110;
   assign mem[409503:409472] = 32'b11111101000101100011000100110100;
   assign mem[409535:409504] = 32'b00000110100111110100010111011000;
   assign mem[409567:409536] = 32'b11111011110000000010111100101000;
   assign mem[409599:409568] = 32'b11111010101101011101101111000000;
   assign mem[409631:409600] = 32'b00000000001001001001110101010101;
   assign mem[409663:409632] = 32'b11111010011110101001110101110000;
   assign mem[409695:409664] = 32'b00000010000001001001111110000100;
   assign mem[409727:409696] = 32'b00000001101110110001001101100110;
   assign mem[409759:409728] = 32'b11111101000001111010000111110000;
   assign mem[409791:409760] = 32'b11111111011011110100111000110110;
   assign mem[409823:409792] = 32'b00000010001100000010100010101100;
   assign mem[409855:409824] = 32'b11111111001000011011000000000101;
   assign mem[409887:409856] = 32'b11111100011011000000110111111000;
   assign mem[409919:409888] = 32'b00000000100010111100001011100000;
   assign mem[409951:409920] = 32'b11111000010111011001000001011000;
   assign mem[409983:409952] = 32'b11111110000101111111111111010110;
   assign mem[410015:409984] = 32'b11111101001110010101111100100100;
   assign mem[410047:410016] = 32'b11111100010000011001011111101100;
   assign mem[410079:410048] = 32'b00000001010111001110111001001010;
   assign mem[410111:410080] = 32'b00000000010011101010100001010110;
   assign mem[410143:410112] = 32'b11111111011111111111110100010110;
   assign mem[410175:410144] = 32'b00001001001100100000100001100000;
   assign mem[410207:410176] = 32'b11111110001001010001000111100000;
   assign mem[410239:410208] = 32'b00000000011000100000100000000001;
   assign mem[410271:410240] = 32'b00000110000011000111011111011000;
   assign mem[410303:410272] = 32'b11110110111011101111010000100000;
   assign mem[410335:410304] = 32'b11111001101000110001100001110000;
   assign mem[410367:410336] = 32'b00000001001001011010100111000010;
   assign mem[410399:410368] = 32'b00000001001011011010100010101110;
   assign mem[410431:410400] = 32'b11111110110100111000001010111010;
   assign mem[410463:410432] = 32'b00000010011010111011010011011000;
   assign mem[410495:410464] = 32'b11110010010010011101011001010000;
   assign mem[410527:410496] = 32'b00001010010101000011011101010000;
   assign mem[410559:410528] = 32'b00000010100001001001000110000100;
   assign mem[410591:410560] = 32'b11111101100001000100110111101100;
   assign mem[410623:410592] = 32'b00001010001110010111100001110000;
   assign mem[410655:410624] = 32'b11111101000011000011001110111000;
   assign mem[410687:410656] = 32'b11111111010000101101010111110111;
   assign mem[410719:410688] = 32'b00000001101011000110010000111010;
   assign mem[410751:410720] = 32'b11111111110001110110110111101010;
   assign mem[410783:410752] = 32'b00000010000011010100110000000000;
   assign mem[410815:410784] = 32'b11111100011111011000100100001000;
   assign mem[410847:410816] = 32'b11111111000011111001111010001000;
   assign mem[410879:410848] = 32'b11111100101010111011000011111000;
   assign mem[410911:410880] = 32'b00000001011001011100011001110110;
   assign mem[410943:410912] = 32'b00000111111011011111000010100000;
   assign mem[410975:410944] = 32'b11111101011000111110101000010100;
   assign mem[411007:410976] = 32'b11111110001001110110011011010010;
   assign mem[411039:411008] = 32'b00000110100001010110011101111000;
   assign mem[411071:411040] = 32'b00000011010111011000110100010100;
   assign mem[411103:411072] = 32'b11111111111100010111011110110001;
   assign mem[411135:411104] = 32'b00000100111100101101001001001000;
   assign mem[411167:411136] = 32'b11110101101110111110001000000000;
   assign mem[411199:411168] = 32'b11111111111001100100011010111000;
   assign mem[411231:411200] = 32'b00010000000011010100101010100000;
   assign mem[411263:411232] = 32'b11111101001100111111000000101100;
   assign mem[411295:411264] = 32'b00000111111101000011011011010000;
   assign mem[411327:411296] = 32'b00000001011010000111011110010000;
   assign mem[411359:411328] = 32'b11110001101111001001010011110000;
   assign mem[411391:411360] = 32'b11111000000000101110010100101000;
   assign mem[411423:411392] = 32'b11111001101011001001110011110000;
   assign mem[411455:411424] = 32'b11111100011110100100001000100100;
   assign mem[411487:411456] = 32'b00000100011001011100000101011000;
   assign mem[411519:411488] = 32'b11110010001110100110110001000000;
   assign mem[411551:411520] = 32'b00000100010101010101101011111000;
   assign mem[411583:411552] = 32'b00001011101000100011101011110000;
   assign mem[411615:411584] = 32'b00000010111000010110100111101000;
   assign mem[411647:411616] = 32'b11111010100001010101011101100000;
   assign mem[411679:411648] = 32'b00000001001010000001010101011100;
   assign mem[411711:411680] = 32'b11110101001100010010000001010000;
   assign mem[411743:411712] = 32'b11111101100010011011000010011100;
   assign mem[411775:411744] = 32'b11111111111001010111101011101111;
   assign mem[411807:411776] = 32'b00000010100010010001010010011100;
   assign mem[411839:411808] = 32'b11111101100000001010010011101000;
   assign mem[411871:411840] = 32'b11110110100101111001101111000000;
   assign mem[411903:411872] = 32'b00001001101011101110001110100000;
   assign mem[411935:411904] = 32'b00000011000010010100101101101000;
   assign mem[411967:411936] = 32'b11110000101010010101111010110000;
   assign mem[411999:411968] = 32'b00000100101001011110011111010000;
   assign mem[412031:412000] = 32'b00000001011010000011100001111110;
   assign mem[412063:412032] = 32'b11111110101010110011100101011010;
   assign mem[412095:412064] = 32'b11111100111010111101111001110100;
   assign mem[412127:412096] = 32'b00000011110011101000110111101000;
   assign mem[412159:412128] = 32'b11111101100001110111111000010100;
   assign mem[412191:412160] = 32'b11110100110100011100110001110000;
   assign mem[412223:412192] = 32'b00001001111110001100111010000000;
   assign mem[412255:412224] = 32'b11101011101110011011110010100000;
   assign mem[412287:412256] = 32'b00001001000110100011010001110000;
   assign mem[412319:412288] = 32'b00000001011100010000101000100100;
   assign mem[412351:412320] = 32'b00000100111101011000000100001000;
   assign mem[412383:412352] = 32'b11111011101101111011111110011000;
   assign mem[412415:412384] = 32'b00000011011110111100010000011100;
   assign mem[412447:412416] = 32'b11110111010000111010000000010000;
   assign mem[412479:412448] = 32'b11111111011010101100110010010110;
   assign mem[412511:412480] = 32'b00000101101011101000000000010000;
   assign mem[412543:412512] = 32'b00000110100101110110111000000000;
   assign mem[412575:412544] = 32'b00000110101000001001001001010000;
   assign mem[412607:412576] = 32'b11111100100011110100110001000000;
   assign mem[412639:412608] = 32'b00000000001010011111010101010100;
   assign mem[412671:412640] = 32'b11111010010010110001010100011000;
   assign mem[412703:412672] = 32'b00000001000111100000001001110110;
   assign mem[412735:412704] = 32'b11111111101001110100000010000011;
   assign mem[412767:412736] = 32'b11111110001011001110000110101110;
   assign mem[412799:412768] = 32'b11111101000110010001010000001100;
   assign mem[412831:412800] = 32'b11111111100011010011001010110100;
   assign mem[412863:412832] = 32'b00001111001101100000001110010000;
   assign mem[412895:412864] = 32'b11111111100000001000100110011111;
   assign mem[412927:412896] = 32'b00000001010011101111100001011100;
   assign mem[412959:412928] = 32'b11111001010110110100100010010000;
   assign mem[412991:412960] = 32'b00000101010100100110110011000000;
   assign mem[413023:412992] = 32'b11111011101100111011111000110000;
   assign mem[413055:413024] = 32'b11111101111010100110001110101100;
   assign mem[413087:413056] = 32'b00000000001110010000010111111000;
   assign mem[413119:413088] = 32'b11111010100011001111101100101000;
   assign mem[413151:413120] = 32'b00000000101001001111111010101100;
   assign mem[413183:413152] = 32'b00000001000011110010011110110100;
   assign mem[413215:413184] = 32'b11111011001101000111101110010000;
   assign mem[413247:413216] = 32'b00000101011101010101101100111000;
   assign mem[413279:413248] = 32'b11111111001011001110011001000100;
   assign mem[413311:413280] = 32'b00000010111010010000101000110100;
   assign mem[413343:413312] = 32'b00000000111110010110000011100101;
   assign mem[413375:413344] = 32'b11111000010000000000001101011000;
   assign mem[413407:413376] = 32'b11111101011001110110010111100100;
   assign mem[413439:413408] = 32'b11111111011011100001001111000000;
   assign mem[413471:413440] = 32'b11111100110101111101110001110100;
   assign mem[413503:413472] = 32'b00000001110011011000001010100100;
   assign mem[413535:413504] = 32'b11110110001011111010011111010000;
   assign mem[413567:413536] = 32'b00010010101011100100101100100000;
   assign mem[413599:413568] = 32'b11110010111000001011011011010000;
   assign mem[413631:413600] = 32'b00000111101111011100101001111000;
   assign mem[413663:413632] = 32'b11110100111010111010001110110000;
   assign mem[413695:413664] = 32'b11110100101001100000000010100000;
   assign mem[413727:413696] = 32'b11111101011011111101000111011000;
   assign mem[413759:413728] = 32'b00000010101101000011001111011000;
   assign mem[413791:413760] = 32'b11110110000101010010011010000000;
   assign mem[413823:413792] = 32'b00000110100010111100111011011000;
   assign mem[413855:413824] = 32'b11100110011110010000101100000000;
   assign mem[413887:413856] = 32'b00010100110000001000001110100000;
   assign mem[413919:413888] = 32'b11111001111100101000100110100000;
   assign mem[413951:413920] = 32'b00000111111000011101110011000000;
   assign mem[413983:413952] = 32'b11111001111000100000000111110000;
   assign mem[414015:413984] = 32'b11111011100011001000111000110000;
   assign mem[414047:414016] = 32'b11101011001100110011111000100000;
   assign mem[414079:414048] = 32'b00000010101001100001011111111100;
   assign mem[414111:414080] = 32'b00000011001001110011101101010000;
   assign mem[414143:414112] = 32'b00000100111111100001000011100000;
   assign mem[414175:414144] = 32'b00000100100000101101110101110000;
   assign mem[414207:414176] = 32'b00000001010100110010110101000100;
   assign mem[414239:414208] = 32'b00000000001111111000011011000000;
   assign mem[414271:414240] = 32'b00000010010100011100110110110100;
   assign mem[414303:414272] = 32'b00000010010011011001110000110000;
   assign mem[414335:414304] = 32'b11111100100110111110010111110000;
   assign mem[414367:414336] = 32'b11111001111010010000000000000000;
   assign mem[414399:414368] = 32'b00000101110011011111100100011000;
   assign mem[414431:414400] = 32'b00000100111000101110011011011000;
   assign mem[414463:414432] = 32'b11111111001101011111110111011000;
   assign mem[414495:414464] = 32'b00000011011000111001000110101000;
   assign mem[414527:414496] = 32'b11111000111101100110011011001000;
   assign mem[414559:414528] = 32'b11110100110010000001100001110000;
   assign mem[414591:414560] = 32'b11111000101111101100000011011000;
   assign mem[414623:414592] = 32'b11111110011111111010000000001010;
   assign mem[414655:414624] = 32'b00000100100001100101000111111000;
   assign mem[414687:414656] = 32'b11111110010001000011000110001000;
   assign mem[414719:414688] = 32'b11111101110010011111101010101100;
   assign mem[414751:414720] = 32'b00000001011101000000110111110010;
   assign mem[414783:414752] = 32'b00000011011101100010111001011100;
   assign mem[414815:414784] = 32'b00000011000000111000101101101000;
   assign mem[414847:414816] = 32'b11111110000101111111001001111100;
   assign mem[414879:414848] = 32'b00000011100101111110000000100100;
   assign mem[414911:414880] = 32'b11111111111001111000010101100010;
   assign mem[414943:414912] = 32'b11111100110110101100110100101100;
   assign mem[414975:414944] = 32'b11111101000001010111010111010100;
   assign mem[415007:414976] = 32'b11111111000101110000101101110110;
   assign mem[415039:415008] = 32'b11111101101110001001100101000100;
   assign mem[415071:415040] = 32'b00000101001000100100100001110000;
   assign mem[415103:415072] = 32'b11110011101000010110101110110000;
   assign mem[415135:415104] = 32'b00000001010101001000100101011110;
   assign mem[415167:415136] = 32'b00000011101101010000000110100000;
   assign mem[415199:415168] = 32'b11110101110110011010111010110000;
   assign mem[415231:415200] = 32'b11111111100010111010110101111000;
   assign mem[415263:415232] = 32'b00000000111011001000010101011100;
   assign mem[415295:415264] = 32'b11111011010011001000100101010000;
   assign mem[415327:415296] = 32'b00000100000101011100100100101000;
   assign mem[415359:415328] = 32'b11111000110010010111111101100000;
   assign mem[415391:415360] = 32'b00000001000001110111101100101010;
   assign mem[415423:415392] = 32'b00000110111110101101111110100000;
   assign mem[415455:415424] = 32'b11111010111001110111010111001000;
   assign mem[415487:415456] = 32'b11111111001111110000001000100000;
   assign mem[415519:415488] = 32'b00000111101110000111010101110000;
   assign mem[415551:415520] = 32'b11111011000001101100000001101000;
   assign mem[415583:415552] = 32'b00000011111001100111011111111100;
   assign mem[415615:415584] = 32'b00000010110000110110011100101100;
   assign mem[415647:415616] = 32'b11110011001100011110111010000000;
   assign mem[415679:415648] = 32'b00000010001100011110001100000100;
   assign mem[415711:415680] = 32'b11111011101110001111101010001000;
   assign mem[415743:415712] = 32'b00000110010111010011101101010000;
   assign mem[415775:415744] = 32'b11111110110110001011011000110000;
   assign mem[415807:415776] = 32'b11111001110110011101000110101000;
   assign mem[415839:415808] = 32'b00000111100100010110000010000000;
   assign mem[415871:415840] = 32'b00000100101011101110001111001000;
   assign mem[415903:415872] = 32'b11110011101000110000111100000000;
   assign mem[415935:415904] = 32'b00001000100001010111001011010000;
   assign mem[415967:415936] = 32'b11110100001001101000111000000000;
   assign mem[415999:415968] = 32'b11111101011101110011001101000000;
   assign mem[416031:416000] = 32'b00000111111101110101101101111000;
   assign mem[416063:416032] = 32'b00000001101110011110110010100000;
   assign mem[416095:416064] = 32'b00000000110010111100011001000101;
   assign mem[416127:416096] = 32'b11111110111101100010111101011010;
   assign mem[416159:416128] = 32'b11110100001010001011101101000000;
   assign mem[416191:416160] = 32'b11111000111111111011101100000000;
   assign mem[416223:416192] = 32'b00000100100110000000011001100000;
   assign mem[416255:416224] = 32'b11111110101110011101101001101110;
   assign mem[416287:416256] = 32'b00000001010100000100110010001110;
   assign mem[416319:416288] = 32'b11111001001001001011011011010000;
   assign mem[416351:416320] = 32'b11111101000110001010110010011000;
   assign mem[416383:416352] = 32'b00001011101100001000100001010000;
   assign mem[416415:416384] = 32'b11110000111100101111111000010000;
   assign mem[416447:416416] = 32'b00000001101010000010100111011010;
   assign mem[416479:416448] = 32'b11111100010010001010001100011100;
   assign mem[416511:416480] = 32'b00000101000111100001101111010000;
   assign mem[416543:416512] = 32'b11110001100101101101111111100000;
   assign mem[416575:416544] = 32'b00000000010101100010111001100111;
   assign mem[416607:416576] = 32'b11111101101010100011011001000000;
   assign mem[416639:416608] = 32'b11111101000011010111011000000100;
   assign mem[416671:416640] = 32'b00000001010010110011110010100110;
   assign mem[416703:416672] = 32'b00000000111100000011100111010011;
   assign mem[416735:416704] = 32'b00001000100110100001111001010000;
   assign mem[416767:416736] = 32'b11111101001100100011010011101000;
   assign mem[416799:416768] = 32'b00000001100100001011011101010100;
   assign mem[416831:416800] = 32'b11111111110001101111010100001010;
   assign mem[416863:416832] = 32'b00000000001000011011111101110000;
   assign mem[416895:416864] = 32'b11111011011110011100110001011000;
   assign mem[416927:416896] = 32'b11111011001100011011011000100000;
   assign mem[416959:416928] = 32'b00000001101000010011000100000100;
   assign mem[416991:416960] = 32'b00000100010111101101101110100000;
   assign mem[417023:416992] = 32'b11101111110111000000001110000000;
   assign mem[417055:417024] = 32'b00001010110001111011001111010000;
   assign mem[417087:417056] = 32'b00000001001000110010101001011110;
   assign mem[417119:417088] = 32'b11111011001001000001010100010000;
   assign mem[417151:417120] = 32'b11111101101000011101101001111000;
   assign mem[417183:417152] = 32'b11111011011011100011000000101000;
   assign mem[417215:417184] = 32'b11110100010101110001101110110000;
   assign mem[417247:417216] = 32'b00000101010010100110000111001000;
   assign mem[417279:417248] = 32'b11111101011001010110101101000000;
   assign mem[417311:417280] = 32'b00000001101000100001001010010000;
   assign mem[417343:417312] = 32'b11110111111110101001001100000000;
   assign mem[417375:417344] = 32'b00000001010110011101111111111000;
   assign mem[417407:417376] = 32'b00000101001001001000010000001000;
   assign mem[417439:417408] = 32'b11110011010001000010101111000000;
   assign mem[417471:417440] = 32'b00000000010000101111000100010111;
   assign mem[417503:417472] = 32'b11111110000101100001101010100110;
   assign mem[417535:417504] = 32'b11101101000110100111001011100000;
   assign mem[417567:417536] = 32'b00000101110100100110110111011000;
   assign mem[417599:417568] = 32'b11111110100010001001011010111110;
   assign mem[417631:417600] = 32'b11111110011011100000001001111000;
   assign mem[417663:417632] = 32'b11111100111101110100111011100100;
   assign mem[417695:417664] = 32'b00001100100011011110011111000000;
   assign mem[417727:417696] = 32'b11101100000001010010110001100000;
   assign mem[417759:417728] = 32'b00000111110001010000101101101000;
   assign mem[417791:417760] = 32'b00000100001000000101000000101000;
   assign mem[417823:417792] = 32'b11111100100001111101111000001000;
   assign mem[417855:417824] = 32'b11111100101101000110010101110000;
   assign mem[417887:417856] = 32'b11111001101000100010000110001000;
   assign mem[417919:417888] = 32'b11111010010000001010100010100000;
   assign mem[417951:417920] = 32'b00000010111110001100100001010100;
   assign mem[417983:417952] = 32'b11111011001111011111110011000000;
   assign mem[418015:417984] = 32'b00001100101111110010110011100000;
   assign mem[418047:418016] = 32'b00000001011000010100001101111110;
   assign mem[418079:418048] = 32'b11111001110000100000010101011000;
   assign mem[418111:418080] = 32'b11110100100011010101101111010000;
   assign mem[418143:418112] = 32'b00000000000001101111100011111011;
   assign mem[418175:418144] = 32'b11101010001001100111101100000000;
   assign mem[418207:418176] = 32'b11111101011000101001000010111100;
   assign mem[418239:418208] = 32'b11110001000011101001110110110000;
   assign mem[418271:418240] = 32'b11101101101111001010001100000000;
   assign mem[418303:418272] = 32'b00000110010111000011111111111000;
   assign mem[418335:418304] = 32'b11111111001111100011110101011000;
   assign mem[418367:418336] = 32'b00000010010110111001011101001000;
   assign mem[418399:418368] = 32'b00000011000001101000011110110000;
   assign mem[418431:418400] = 32'b00000110111010110010001110000000;
   assign mem[418463:418432] = 32'b11101110010010111101100010000000;
   assign mem[418495:418464] = 32'b00000011101111101110011000000000;
   assign mem[418527:418496] = 32'b00000001110101011110100000101100;
   assign mem[418559:418528] = 32'b00000100101100111100010010101000;
   assign mem[418591:418560] = 32'b00000011101100000110101001110100;
   assign mem[418623:418592] = 32'b00000011001100010000010100010100;
   assign mem[418655:418624] = 32'b00000011110000010001011111101100;
   assign mem[418687:418656] = 32'b11111110010001100000010001010000;
   assign mem[418719:418688] = 32'b11111110011000111010011111100000;
   assign mem[418751:418720] = 32'b11111110111010101000100011100000;
   assign mem[418783:418752] = 32'b00000001010100111001000101011000;
   assign mem[418815:418784] = 32'b11111110011110110101010000001110;
   assign mem[418847:418816] = 32'b11111001011010010001001011001000;
   assign mem[418879:418848] = 32'b11111101111000001001010000101000;
   assign mem[418911:418880] = 32'b11111000010100110100110001010000;
   assign mem[418943:418912] = 32'b00000101101100010000110110010000;
   assign mem[418975:418944] = 32'b11110100101010101100101010010000;
   assign mem[419007:418976] = 32'b00001101000010001011101010000000;
   assign mem[419039:419008] = 32'b11111001110001000101010101001000;
   assign mem[419071:419040] = 32'b00000010001101100101000000111000;
   assign mem[419103:419072] = 32'b11101010111110101001111111100000;
   assign mem[419135:419104] = 32'b11111011010110000010111101110000;
   assign mem[419167:419136] = 32'b11110001000000011100011111010000;
   assign mem[419199:419168] = 32'b00000101010010100011101000100000;
   assign mem[419231:419200] = 32'b00001001010100010000011100000000;
   assign mem[419263:419232] = 32'b11111010011110001111011101010000;
   assign mem[419295:419264] = 32'b11111111110000001010010101100010;
   assign mem[419327:419296] = 32'b11111000011101110000100110010000;
   assign mem[419359:419328] = 32'b11111010111111011010001001110000;
   assign mem[419391:419360] = 32'b11111001100100111101000010100000;
   assign mem[419423:419392] = 32'b11110111111010000001111001000000;
   assign mem[419455:419424] = 32'b00000000101001000011010111001001;
   assign mem[419487:419456] = 32'b11111111100011000011101101010101;
   assign mem[419519:419488] = 32'b00000010001000011001011010001000;
   assign mem[419551:419520] = 32'b11111111110010100011101011100101;
   assign mem[419583:419552] = 32'b00000100110011011000111011111000;
   assign mem[419615:419584] = 32'b11111111101010100000101001011100;
   assign mem[419647:419616] = 32'b11111111010001101101010110010010;
   assign mem[419679:419648] = 32'b11111110111001100011001011110000;
   assign mem[419711:419680] = 32'b11111110011101101010100110101110;
   assign mem[419743:419712] = 32'b11111010111101000011010111010000;
   assign mem[419775:419744] = 32'b11110111000110110110101000010000;
   assign mem[419807:419776] = 32'b00000011100111000010100111110000;
   assign mem[419839:419808] = 32'b00000000001100000100101100010000;
   assign mem[419871:419840] = 32'b00000100011010011101011011001000;
   assign mem[419903:419872] = 32'b00001010110011100011110011110000;
   assign mem[419935:419904] = 32'b00000001110010100110011100111100;
   assign mem[419967:419936] = 32'b11110111010111011011010111010000;
   assign mem[419999:419968] = 32'b00000100000011001101110010101000;
   assign mem[420031:420000] = 32'b00000011001010111110101100110000;
   assign mem[420063:420032] = 32'b11110100001100101011111001010000;
   assign mem[420095:420064] = 32'b00000100010011111100011101111000;
   assign mem[420127:420096] = 32'b00000100111110001101010010001000;
   assign mem[420159:420128] = 32'b11110100111000100001011111100000;
   assign mem[420191:420160] = 32'b00001100000101001000000010010000;
   assign mem[420223:420192] = 32'b00000010100110001101110100101000;
   assign mem[420255:420224] = 32'b00000001100110100000001010100110;
   assign mem[420287:420256] = 32'b11110110111010111100000010100000;
   assign mem[420319:420288] = 32'b11110110110110110011101000000000;
   assign mem[420351:420320] = 32'b11110100101111110110011001010000;
   assign mem[420383:420352] = 32'b11111110000001101001101100001100;
   assign mem[420415:420384] = 32'b00001010001110110111111000010000;
   assign mem[420447:420416] = 32'b11111110001001001101010000000100;
   assign mem[420479:420448] = 32'b11111101011001110110110110100100;
   assign mem[420511:420480] = 32'b00000011011011010001010110011100;
   assign mem[420543:420512] = 32'b00000111000100110001011101001000;
   assign mem[420575:420544] = 32'b00000000001100111011110011010111;
   assign mem[420607:420576] = 32'b11111111101001110101101000010100;
   assign mem[420639:420608] = 32'b11111110111110001010001001101110;
   assign mem[420671:420640] = 32'b00000011011001110001000010001000;
   assign mem[420703:420672] = 32'b00000001011010001100111111011100;
   assign mem[420735:420704] = 32'b11111010000110101111110101110000;
   assign mem[420767:420736] = 32'b00000010000011111000000110001100;
   assign mem[420799:420768] = 32'b00000000100110100000101100100101;
   assign mem[420831:420800] = 32'b11110000010110100100101100000000;
   assign mem[420863:420832] = 32'b00000101101000011001000011001000;
   assign mem[420895:420864] = 32'b00000100110110110100100111100000;
   assign mem[420927:420896] = 32'b11111001010100110011110000110000;
   assign mem[420959:420928] = 32'b00000010110010010011000010000100;
   assign mem[420991:420960] = 32'b00000101101011000100111000000000;
   assign mem[421023:420992] = 32'b11101111001010100100100001000000;
   assign mem[421055:421024] = 32'b11111111010011110111111101101101;
   assign mem[421087:421056] = 32'b11111010011100010000110001000000;
   assign mem[421119:421088] = 32'b00000001000110001000100100100010;
   assign mem[421151:421120] = 32'b00000001101000110011010110101110;
   assign mem[421183:421152] = 32'b00000011001111000100111110010000;
   assign mem[421215:421184] = 32'b11111110110110011110111111111110;
   assign mem[421247:421216] = 32'b00000100010110000110001011101000;
   assign mem[421279:421248] = 32'b11111111101000001101001101100101;
   assign mem[421311:421280] = 32'b00000011011111000010101001000000;
   assign mem[421343:421312] = 32'b11111011011011000101101001100000;
   assign mem[421375:421344] = 32'b00000000010001001011101000001010;
   assign mem[421407:421376] = 32'b11110000100000101010011000100000;
   assign mem[421439:421408] = 32'b11111110001011001000111110000000;
   assign mem[421471:421440] = 32'b11110101011010110011010111100000;
   assign mem[421503:421472] = 32'b00000111101110010101101010111000;
   assign mem[421535:421504] = 32'b11111110001100011111110100111010;
   assign mem[421567:421536] = 32'b00000011100110111001001110011000;
   assign mem[421599:421568] = 32'b00000000100001110011010110110100;
   assign mem[421631:421600] = 32'b00000011110101110101000100111100;
   assign mem[421663:421632] = 32'b11110101011010101110101000010000;
   assign mem[421695:421664] = 32'b11111001000101101001001001101000;
   assign mem[421727:421696] = 32'b11111010000000110111000001100000;
   assign mem[421759:421728] = 32'b00000111100010010100010001011000;
   assign mem[421791:421760] = 32'b11111110110101110110100111100100;
   assign mem[421823:421792] = 32'b11111101101000011100001011110100;
   assign mem[421855:421824] = 32'b00000010010100101100110001101000;
   assign mem[421887:421856] = 32'b00000111001011011001101011101000;
   assign mem[421919:421888] = 32'b00000110110001111101001011010000;
   assign mem[421951:421920] = 32'b00000000001110000101100001101011;
   assign mem[421983:421952] = 32'b11111011110101011101011010101000;
   assign mem[422015:421984] = 32'b11110110101100101011010001000000;
   assign mem[422047:422016] = 32'b11110111100101110000010101110000;
   assign mem[422079:422048] = 32'b11111101111011100110100011011100;
   assign mem[422111:422080] = 32'b11111101010010111111011000101000;
   assign mem[422143:422112] = 32'b00001000100100011000010010000000;
   assign mem[422175:422144] = 32'b11111100100000100010001000111100;
   assign mem[422207:422176] = 32'b00000111111001111010101101101000;
   assign mem[422239:422208] = 32'b00000100001001010101111101010000;
   assign mem[422271:422240] = 32'b11111111111100001001111110110101;
   assign mem[422303:422272] = 32'b11110101100110001101011010010000;
   assign mem[422335:422304] = 32'b00000011001001111101110001110000;
   assign mem[422367:422336] = 32'b11110100001000101010011010000000;
   assign mem[422399:422368] = 32'b00000000010000100001001111100101;
   assign mem[422431:422400] = 32'b00000000110110110100000010000111;
   assign mem[422463:422432] = 32'b11101100011010110101010010100000;
   assign mem[422495:422464] = 32'b00000001001100011000000001000000;
   assign mem[422527:422496] = 32'b00000010010011111001100110110100;
   assign mem[422559:422528] = 32'b00000000010001000000100101010110;
   assign mem[422591:422560] = 32'b11111110110010101010000100100010;
   assign mem[422623:422592] = 32'b00000000110001100011010111101111;
   assign mem[422655:422624] = 32'b11110010100101111011011001000000;
   assign mem[422687:422656] = 32'b00000100011111100010100001011000;
   assign mem[422719:422688] = 32'b11111110111111110011000110100000;
   assign mem[422751:422720] = 32'b00000010011010110110101101101000;
   assign mem[422783:422752] = 32'b00000110100101011111000110110000;
   assign mem[422815:422784] = 32'b11111110011101010000100101010000;
   assign mem[422847:422816] = 32'b11111101011000111100101111010100;
   assign mem[422879:422848] = 32'b00000001101110011111110010101110;
   assign mem[422911:422880] = 32'b00000100011010000101011001010000;
   assign mem[422943:422912] = 32'b00000010010000011000110101100000;
   assign mem[422975:422944] = 32'b11111010110011010010011010100000;
   assign mem[423007:422976] = 32'b11111000000111100101110111001000;
   assign mem[423039:423008] = 32'b11111101110111100001101100110100;
   assign mem[423071:423040] = 32'b00000001001101110010101110001100;
   assign mem[423103:423072] = 32'b00000010100110001101010111000100;
   assign mem[423135:423104] = 32'b00000000000100000010001100111100;
   assign mem[423167:423136] = 32'b11111101010100111001001000011100;
   assign mem[423199:423168] = 32'b00000010101011100110111011010000;
   assign mem[423231:423200] = 32'b11111111011101111010000010111101;
   assign mem[423263:423232] = 32'b11111111011100110100111010101001;
   assign mem[423295:423264] = 32'b11111011001000010101100111101000;
   assign mem[423327:423296] = 32'b00000010111010011110110000111100;
   assign mem[423359:423328] = 32'b00000000011011001000010110101000;
   assign mem[423391:423360] = 32'b11111110100011000111000000110000;
   assign mem[423423:423392] = 32'b00000101100000011100101000010000;
   assign mem[423455:423424] = 32'b00000110011110010100101001010000;
   assign mem[423487:423456] = 32'b00000110100001110100010010010000;
   assign mem[423519:423488] = 32'b00000011111101100010000010011000;
   assign mem[423551:423520] = 32'b11110011111101000100100010010000;
   assign mem[423583:423552] = 32'b00000011010001110010001100000000;
   assign mem[423615:423584] = 32'b11111011100001111101100010101000;
   assign mem[423647:423616] = 32'b11111101100111011011000011001000;
   assign mem[423679:423648] = 32'b11111111011110011010100101111111;
   assign mem[423711:423680] = 32'b00000001101011110101100110101000;
   assign mem[423743:423712] = 32'b11110001100100001111010100000000;
   assign mem[423775:423744] = 32'b11111110000011101011001110001100;
   assign mem[423807:423776] = 32'b00000000000010100011100100001100;
   assign mem[423839:423808] = 32'b11111110110100111101100101111010;
   assign mem[423871:423840] = 32'b00000000100110001001010010001011;
   assign mem[423903:423872] = 32'b00000000100010011011000111001010;
   assign mem[423935:423904] = 32'b11111100100001100011000100010000;
   assign mem[423967:423936] = 32'b00000100110000011010011010001000;
   assign mem[423999:423968] = 32'b00000000010011010010000110001010;
   assign mem[424031:424000] = 32'b11111101100101110000001101110100;
   assign mem[424063:424032] = 32'b00000001101001110001011101100110;
   assign mem[424095:424064] = 32'b00000000000101101111110001100111;
   assign mem[424127:424096] = 32'b00000001111101100110100001000100;
   assign mem[424159:424128] = 32'b11111010100111001111101100001000;
   assign mem[424191:424160] = 32'b00000100010011000111001100110000;
   assign mem[424223:424192] = 32'b11110111011000101000100101010000;
   assign mem[424255:424224] = 32'b00000100011000011101011000101000;
   assign mem[424287:424256] = 32'b00000000101011001101010010001110;
   assign mem[424319:424288] = 32'b11111001101111010101111010011000;
   assign mem[424351:424320] = 32'b00000110101100110110111101000000;
   assign mem[424383:424352] = 32'b00000001110110010101101001111110;
   assign mem[424415:424384] = 32'b00000111011111101000010100001000;
   assign mem[424447:424416] = 32'b00000110011110100011000101101000;
   assign mem[424479:424448] = 32'b11111110010000011111001110100100;
   assign mem[424511:424480] = 32'b11111101000000010001110100011100;
   assign mem[424543:424512] = 32'b00000010010100110010111100111000;
   assign mem[424575:424544] = 32'b11110010111011011000010001000000;
   assign mem[424607:424576] = 32'b00000001110000011111000111010110;
   assign mem[424639:424608] = 32'b11111000011000001011111110000000;
   assign mem[424671:424640] = 32'b11111111000101000101100001101010;
   assign mem[424703:424672] = 32'b11111110011010010010111011111000;
   assign mem[424735:424704] = 32'b00000001001111110111111011101100;
   assign mem[424767:424736] = 32'b11111110100100110011111100010000;
   assign mem[424799:424768] = 32'b11111101100110000111001001000000;
   assign mem[424831:424800] = 32'b00000001100110100010100001001010;
   assign mem[424863:424832] = 32'b00000000001001011011011111010001;
   assign mem[424895:424864] = 32'b00000011011011001000011101100100;
   assign mem[424927:424896] = 32'b11111110000011001110011001001100;
   assign mem[424959:424928] = 32'b11111100100100010000111110001100;
   assign mem[424991:424960] = 32'b00000010000011101011111110101000;
   assign mem[425023:424992] = 32'b11111001010101111001010101110000;
   assign mem[425055:425024] = 32'b00001000010011110100100100100000;
   assign mem[425087:425056] = 32'b11111000010010111110000111111000;
   assign mem[425119:425088] = 32'b00001000010011111100010001010000;
   assign mem[425151:425120] = 32'b11111100100100000001100100011100;
   assign mem[425183:425152] = 32'b00000000011001000100011110000011;
   assign mem[425215:425184] = 32'b11111100000111011100101110111000;
   assign mem[425247:425216] = 32'b11111001000111011101011010011000;
   assign mem[425279:425248] = 32'b11111110000111111110101000000000;
   assign mem[425311:425280] = 32'b11111001100111000011010010000000;
   assign mem[425343:425312] = 32'b00000011011010011010101010110000;
   assign mem[425375:425344] = 32'b00000011101011111011011111011100;
   assign mem[425407:425376] = 32'b11111010110000011001110001011000;
   assign mem[425439:425408] = 32'b11110011101111010011010010010000;
   assign mem[425471:425440] = 32'b11110111100101100001001000110000;
   assign mem[425503:425472] = 32'b11111100000000111010011100001000;
   assign mem[425535:425504] = 32'b00001001111010100001001001100000;
   assign mem[425567:425536] = 32'b00000000000011011110110000100110;
   assign mem[425599:425568] = 32'b00000011100001111000111011111000;
   assign mem[425631:425600] = 32'b00000011111111101101101001010100;
   assign mem[425663:425632] = 32'b00000000111010101111101111001010;
   assign mem[425695:425664] = 32'b11111110111111100100101000101000;
   assign mem[425727:425696] = 32'b11110111101010001001001101110000;
   assign mem[425759:425728] = 32'b11111011111011110111011001001000;
   assign mem[425791:425760] = 32'b11111110011000101000001011101110;
   assign mem[425823:425792] = 32'b11111110111100000111001111011010;
   assign mem[425855:425824] = 32'b00000010111010101010001110110000;
   assign mem[425887:425856] = 32'b11111011110001100001001110000000;
   assign mem[425919:425888] = 32'b00000010011110110101110111000100;
   assign mem[425951:425920] = 32'b00000010101100001010000100101100;
   assign mem[425983:425952] = 32'b00000010010011100001110101010000;
   assign mem[426015:425984] = 32'b00000000100001100001110110110111;
   assign mem[426047:426016] = 32'b11111111010100111100001101100100;
   assign mem[426079:426048] = 32'b11111101010101101110000010000000;
   assign mem[426111:426080] = 32'b11111111101010101110111111101010;
   assign mem[426143:426112] = 32'b11111111110100100100010110001001;
   assign mem[426175:426144] = 32'b11110111010101100000011101000000;
   assign mem[426207:426176] = 32'b00000001001111001100010001011100;
   assign mem[426239:426208] = 32'b11111111001011100011110101011010;
   assign mem[426271:426240] = 32'b00000001101011000001010101110010;
   assign mem[426303:426272] = 32'b00000000000011011000000101010111;
   assign mem[426335:426304] = 32'b00000100000111010100001000101000;
   assign mem[426367:426336] = 32'b00000000000001010110100100100101;
   assign mem[426399:426368] = 32'b00000000000010000100001100000111;
   assign mem[426431:426400] = 32'b11111011011010001110111110011000;
   assign mem[426463:426432] = 32'b11111010101011010010110000110000;
   assign mem[426495:426464] = 32'b11110110010001110011100111100000;
   assign mem[426527:426496] = 32'b00000010010011100110110001011100;
   assign mem[426559:426528] = 32'b11111100001111100110010110100100;
   assign mem[426591:426560] = 32'b11111101110110010001001011011000;
   assign mem[426623:426592] = 32'b00001010010000010010001011010000;
   assign mem[426655:426624] = 32'b11111011010111011000110111011000;
   assign mem[426687:426656] = 32'b11111111101011010001110000100100;
   assign mem[426719:426688] = 32'b00000011001001010100010011111000;
   assign mem[426751:426720] = 32'b11111110101101101010111110010000;
   assign mem[426783:426752] = 32'b11111111001000110001000000000011;
   assign mem[426815:426784] = 32'b11111100101100000010011000101100;
   assign mem[426847:426816] = 32'b00000010101000110101010000100000;
   assign mem[426879:426848] = 32'b00000001000110110110010101011100;
   assign mem[426911:426880] = 32'b00000010111111110010111111100000;
   assign mem[426943:426912] = 32'b00000010001101001011001101100000;
   assign mem[426975:426944] = 32'b00000010001000101001001101000000;
   assign mem[427007:426976] = 32'b00000000011001001011111010100011;
   assign mem[427039:427008] = 32'b11111110110011110001011000011010;
   assign mem[427071:427040] = 32'b11111100110001100010010111100000;
   assign mem[427103:427072] = 32'b11111110101101011000101101101000;
   assign mem[427135:427104] = 32'b11110111010101011001011001110000;
   assign mem[427167:427136] = 32'b00000110011001110110101101011000;
   assign mem[427199:427168] = 32'b11111001010101110101100101111000;
   assign mem[427231:427200] = 32'b11110110011100001001101101110000;
   assign mem[427263:427232] = 32'b00010001111001011111111000100000;
   assign mem[427295:427264] = 32'b00001001100111001001011111110000;
   assign mem[427327:427296] = 32'b11111101111100111111010100010100;
   assign mem[427359:427328] = 32'b00000011100001001111010000100100;
   assign mem[427391:427360] = 32'b11111010110010100010110011000000;
   assign mem[427423:427392] = 32'b11110000010101001000111111100000;
   assign mem[427455:427424] = 32'b11111101000101000110100111100000;
   assign mem[427487:427456] = 32'b00000001001010010000000011110110;
   assign mem[427519:427488] = 32'b11110111011001010001111011100000;
   assign mem[427551:427520] = 32'b00000010000101011100011100001100;
   assign mem[427583:427552] = 32'b00000001100100101110101100001110;
   assign mem[427615:427584] = 32'b00000011010011111111001111011100;
   assign mem[427647:427616] = 32'b00000100011111000001001000010000;
   assign mem[427679:427648] = 32'b11111010010010001011010010111000;
   assign mem[427711:427680] = 32'b00000000100101101100000100100011;
   assign mem[427743:427712] = 32'b11111110111011110000001101111000;
   assign mem[427775:427744] = 32'b00000000100100111110001001001001;
   assign mem[427807:427776] = 32'b11111011010111000100101000111000;
   assign mem[427839:427808] = 32'b00000000111111001001011111010100;
   assign mem[427871:427840] = 32'b00000001100101010101110110000000;
   assign mem[427903:427872] = 32'b11111101000100011011000111100100;
   assign mem[427935:427904] = 32'b00000001001110011101101101001010;
   assign mem[427967:427936] = 32'b00000010011110001100010101001000;
   assign mem[427999:427968] = 32'b11111011011011010011001001101000;
   assign mem[428031:428000] = 32'b11111111101000011101110001111000;
   assign mem[428063:428032] = 32'b11111110110100001100011100001000;
   assign mem[428095:428064] = 32'b11110010001010100000111111010000;
   assign mem[428127:428096] = 32'b11111111001010011110001011110001;
   assign mem[428159:428128] = 32'b11111111110110011011111101011111;
   assign mem[428191:428160] = 32'b11110000101001001111110000000000;
   assign mem[428223:428192] = 32'b00000100000101011100100110101000;
   assign mem[428255:428224] = 32'b11110001000110010101011010010000;
   assign mem[428287:428256] = 32'b00001010100101110111111101000000;
   assign mem[428319:428288] = 32'b11110111010000101101100101010000;
   assign mem[428351:428320] = 32'b00001000111001101000011001000000;
   assign mem[428383:428352] = 32'b11110011000111101111001010010000;
   assign mem[428415:428384] = 32'b00000010010000011111101110001000;
   assign mem[428447:428416] = 32'b11110000000110011000111110010000;
   assign mem[428479:428448] = 32'b00000101111010100010001000001000;
   assign mem[428511:428480] = 32'b11111001000001001111000100110000;
   assign mem[428543:428512] = 32'b11111111100010110011001001001100;
   assign mem[428575:428544] = 32'b11111100000101100110100011010000;
   assign mem[428607:428576] = 32'b00000100111011001111111110000000;
   assign mem[428639:428608] = 32'b11111110011101011100100110001110;
   assign mem[428671:428640] = 32'b00000001101010110001111011111010;
   assign mem[428703:428672] = 32'b11110001101100011101101100000000;
   assign mem[428735:428704] = 32'b00000001011011010111011100011100;
   assign mem[428767:428736] = 32'b00000000111101110111010001011000;
   assign mem[428799:428768] = 32'b00000110111101010110011111010000;
   assign mem[428831:428800] = 32'b11100001000101111100001001000000;
   assign mem[428863:428832] = 32'b00000101101000001101111100110000;
   assign mem[428895:428864] = 32'b11111010110010100010001110010000;
   assign mem[428927:428896] = 32'b00000011110110101111000011111100;
   assign mem[428959:428928] = 32'b11111111011001100101111101101011;
   assign mem[428991:428960] = 32'b00000101100100101000111011101000;
   assign mem[429023:428992] = 32'b11101000010100101000010111000000;
   assign mem[429055:429024] = 32'b00000001001110101101000101111110;
   assign mem[429087:429056] = 32'b11111011010001000010011010110000;
   assign mem[429119:429088] = 32'b00000101010101101111111111100000;
   assign mem[429151:429120] = 32'b00000011011110111011111001001000;
   assign mem[429183:429152] = 32'b00000000010100011000111111110011;
   assign mem[429215:429184] = 32'b00000010001000010100110001011000;
   assign mem[429247:429216] = 32'b11101111011110110111101101000000;
   assign mem[429279:429248] = 32'b11111111010111000010101110010100;
   assign mem[429311:429280] = 32'b11110100110000101010010010110000;
   assign mem[429343:429312] = 32'b11110111111100001000010000000000;
   assign mem[429375:429344] = 32'b00001000001010101111011000000000;
   assign mem[429407:429376] = 32'b00000011011001000110001110110000;
   assign mem[429439:429408] = 32'b11111111000101111101011010011101;
   assign mem[429471:429440] = 32'b00000111010100100100100010110000;
   assign mem[429503:429472] = 32'b00000010100011010100000011000100;
   assign mem[429535:429504] = 32'b00000110100001011010010011001000;
   assign mem[429567:429536] = 32'b00000010101100111000110000001000;
   assign mem[429599:429568] = 32'b11111000100010001011011111011000;
   assign mem[429631:429600] = 32'b11111011010000010011101111111000;
   assign mem[429663:429632] = 32'b11111111011111000000000101011110;
   assign mem[429695:429664] = 32'b00000000010101110011111001100010;
   assign mem[429727:429696] = 32'b11111111100011100100101000000011;
   assign mem[429759:429728] = 32'b11111011000001100111100000110000;
   assign mem[429791:429760] = 32'b00000010000111001010110101000000;
   assign mem[429823:429792] = 32'b00001011010001011100001011000000;
   assign mem[429855:429824] = 32'b00000101001000100011000001000000;
   assign mem[429887:429856] = 32'b11111101010101101011001011100000;
   assign mem[429919:429888] = 32'b11110111110000001110000000100000;
   assign mem[429951:429920] = 32'b11111001000111101111011000100000;
   assign mem[429983:429952] = 32'b11111110011110100011100100100110;
   assign mem[430015:429984] = 32'b11111010110011011010100000000000;
   assign mem[430047:430016] = 32'b00000000001101100100011000101000;
   assign mem[430079:430048] = 32'b11111100101111101100000100010100;
   assign mem[430111:430080] = 32'b00000001001011111100110100101010;
   assign mem[430143:430112] = 32'b11111011100001111101111001011000;
   assign mem[430175:430144] = 32'b11111110101001100011100101001010;
   assign mem[430207:430176] = 32'b00000010010001101011010110111000;
   assign mem[430239:430208] = 32'b11111101011111111011011010110000;
   assign mem[430271:430240] = 32'b11111111001101110010101111111100;
   assign mem[430303:430272] = 32'b11111110000111001100010010111100;
   assign mem[430335:430304] = 32'b11110110001111010111000000110000;
   assign mem[430367:430336] = 32'b00000011100001110001111010011100;
   assign mem[430399:430368] = 32'b11111101001001100000010101100000;
   assign mem[430431:430400] = 32'b00001011011011001110011100100000;
   assign mem[430463:430432] = 32'b11111100001011001001100001001000;
   assign mem[430495:430464] = 32'b11110101001001011111011101100000;
   assign mem[430527:430496] = 32'b00000010111010001011000110000000;
   assign mem[430559:430528] = 32'b11110100011110011101100111010000;
   assign mem[430591:430560] = 32'b00000010011101001000010010000100;
   assign mem[430623:430592] = 32'b11111110001001110101001010011000;
   assign mem[430655:430624] = 32'b00000101000100001001011100010000;
   assign mem[430687:430656] = 32'b11110101001011110100000100000000;
   assign mem[430719:430688] = 32'b00000110000011111001001100001000;
   assign mem[430751:430720] = 32'b11111110010010110010000000000010;
   assign mem[430783:430752] = 32'b11110101101011101111011011000000;
   assign mem[430815:430784] = 32'b00000011001100001100011011101100;
   assign mem[430847:430816] = 32'b00000010111001011101001001111000;
   assign mem[430879:430848] = 32'b11111111100010001010100110000101;
   assign mem[430911:430880] = 32'b00000010101000100001011110110100;
   assign mem[430943:430912] = 32'b00000100100110000111101101111000;
   assign mem[430975:430944] = 32'b11100010110001111011001111000000;
   assign mem[431007:430976] = 32'b00000110011000011110011101011000;
   assign mem[431039:431008] = 32'b11111101001110010000100100111100;
   assign mem[431071:431040] = 32'b00000000110110101010101010111001;
   assign mem[431103:431072] = 32'b11111101100101010101011100110000;
   assign mem[431135:431104] = 32'b11111100101001101001010100110000;
   assign mem[431167:431136] = 32'b00000010001001100001011100101000;
   assign mem[431199:431168] = 32'b11111100001111010101011000110100;
   assign mem[431231:431200] = 32'b00000100010010010011001000010000;
   assign mem[431263:431232] = 32'b00000001110000010010100000000110;
   assign mem[431295:431264] = 32'b00000000101111100111101000111011;
   assign mem[431327:431296] = 32'b11111011111100100000101011010000;
   assign mem[431359:431328] = 32'b00000100110000001111000110110000;
   assign mem[431391:431360] = 32'b11111111000101001001000100000110;
   assign mem[431423:431392] = 32'b00000000110110000001001010111110;
   assign mem[431455:431424] = 32'b00000010101011011001001111110000;
   assign mem[431487:431456] = 32'b11111111011101110001001000100000;
   assign mem[431519:431488] = 32'b11111110110000000111111101111110;
   assign mem[431551:431520] = 32'b00000011111010010111000001000000;
   assign mem[431583:431552] = 32'b11111100000011011100111011111100;
   assign mem[431615:431584] = 32'b00000000011111011110111110110101;
   assign mem[431647:431616] = 32'b11110111001100111001001111010000;
   assign mem[431679:431648] = 32'b00000101010001111000100000001000;
   assign mem[431711:431680] = 32'b00000000011011010000111010100110;
   assign mem[431743:431712] = 32'b11111110111010100110011111100010;
   assign mem[431775:431744] = 32'b11111111011001111100101011010111;
   assign mem[431807:431776] = 32'b11110101110101010001011000010000;
   assign mem[431839:431808] = 32'b00000100001000001100110011100000;
   assign mem[431871:431840] = 32'b11110111111110011010001011110000;
   assign mem[431903:431872] = 32'b11111010111110011000011010101000;
   assign mem[431935:431904] = 32'b00000110111010101010000001011000;
   assign mem[431967:431936] = 32'b00000011101011000111111111101000;
   assign mem[431999:431968] = 32'b00000000010010111011010010010101;
   assign mem[432031:432000] = 32'b11101111101110001011000011100000;
   assign mem[432063:432032] = 32'b00001111000011111100000000110000;
   assign mem[432095:432064] = 32'b00001010110011001110010101100000;
   assign mem[432127:432096] = 32'b11110011110111010110100011110000;
   assign mem[432159:432128] = 32'b11111110000100001010100011001100;
   assign mem[432191:432160] = 32'b00000000011000000111111000001110;
   assign mem[432223:432192] = 32'b11100110000110101100101111000000;
   assign mem[432255:432224] = 32'b00001101100110000101011011010000;
   assign mem[432287:432256] = 32'b11111101001001110001011010100000;
   assign mem[432319:432288] = 32'b11111010000011010101000101101000;
   assign mem[432351:432320] = 32'b11110110011011011111101111100000;
   assign mem[432383:432352] = 32'b00000101110000110111110001101000;
   assign mem[432415:432384] = 32'b11111100110111010101111110101000;
   assign mem[432447:432416] = 32'b11110111100010000100111000000000;
   assign mem[432479:432448] = 32'b00000010001001111100001010100000;
   assign mem[432511:432480] = 32'b11111100110101011110111110110000;
   assign mem[432543:432512] = 32'b11111001111100110101000101000000;
   assign mem[432575:432544] = 32'b00000101011111000110000001110000;
   assign mem[432607:432576] = 32'b11110110000100111111010000010000;
   assign mem[432639:432608] = 32'b00000011101101011101110110100100;
   assign mem[432671:432640] = 32'b11111110000101000111101111111100;
   assign mem[432703:432672] = 32'b00000110111111000111001111011000;
   assign mem[432735:432704] = 32'b11101100101010100110010111000000;
   assign mem[432767:432736] = 32'b00001001000011011100010111000000;
   assign mem[432799:432768] = 32'b11110101000101101100001001000000;
   assign mem[432831:432800] = 32'b00001001111001110110101111100000;
   assign mem[432863:432832] = 32'b11110010100000001101011100110000;
   assign mem[432895:432864] = 32'b11110101110001111100001100100000;
   assign mem[432927:432896] = 32'b11110000001110111011011000110000;
   assign mem[432959:432928] = 32'b00000011011111000100111001001000;
   assign mem[432991:432960] = 32'b11111111010110101110011011000001;
   assign mem[433023:432992] = 32'b00000101001010100111001100111000;
   assign mem[433055:433024] = 32'b00000101101010010000000110100000;
   assign mem[433087:433056] = 32'b11110000100010001010000000100000;
   assign mem[433119:433088] = 32'b00000000000001010100100111101000;
   assign mem[433151:433120] = 32'b11101100111101010010100100000000;
   assign mem[433183:433152] = 32'b11111001010101001001011101110000;
   assign mem[433215:433184] = 32'b00000001011100110110001001110110;
   assign mem[433247:433216] = 32'b00000011000011011010110110011000;
   assign mem[433279:433248] = 32'b11111110100010111010101110010100;
   assign mem[433311:433280] = 32'b00000010000101111101100100100000;
   assign mem[433343:433312] = 32'b00001001001101110100111100010000;
   assign mem[433375:433344] = 32'b11111001100001100001101010111000;
   assign mem[433407:433376] = 32'b11111111111011010000100010000011;
   assign mem[433439:433408] = 32'b00000010001100110110100111001000;
   assign mem[433471:433440] = 32'b00001000100100110011110110000000;
   assign mem[433503:433472] = 32'b11111001000010011110011010111000;
   assign mem[433535:433504] = 32'b11111001100001000000000110000000;
   assign mem[433567:433536] = 32'b11111100011000100101100010110100;
   assign mem[433599:433568] = 32'b00000011111000001000110111010000;
   assign mem[433631:433600] = 32'b11111110110101010011001011010010;
   assign mem[433663:433632] = 32'b11111100011100011011101001010100;
   assign mem[433695:433664] = 32'b11111101010001001001111001001000;
   assign mem[433727:433696] = 32'b11111110100101101010010111011110;
   assign mem[433759:433728] = 32'b11111001101011001011100011010000;
   assign mem[433791:433760] = 32'b00000001101001110111100101111100;
   assign mem[433823:433792] = 32'b00000011100111010011101000010100;
   assign mem[433855:433824] = 32'b11111000000101100110010110011000;
   assign mem[433887:433856] = 32'b00000000010110010101010001110101;
   assign mem[433919:433888] = 32'b11111110101101011111101011010010;
   assign mem[433951:433920] = 32'b00000111000000100101000000110000;
   assign mem[433983:433952] = 32'b00000011011110001111000010011000;
   assign mem[434015:433984] = 32'b11111110011000000101011011000110;
   assign mem[434047:434016] = 32'b00000000110011101010110110100111;
   assign mem[434079:434048] = 32'b11111000000110001110001111001000;
   assign mem[434111:434080] = 32'b11111111110101001010010111110100;
   assign mem[434143:434112] = 32'b00000010110101010101011010101100;
   assign mem[434175:434144] = 32'b11100111010100001101011001100000;
   assign mem[434207:434176] = 32'b00000110111000100011010111100000;
   assign mem[434239:434208] = 32'b11111100010011100111101011010100;
   assign mem[434271:434240] = 32'b11111010110001100010010110001000;
   assign mem[434303:434272] = 32'b00001100111101111010101000000000;
   assign mem[434335:434304] = 32'b11110111101011111010010001110000;
   assign mem[434367:434336] = 32'b00000100000011100110110100000000;
   assign mem[434399:434368] = 32'b11110001111101001000011011100000;
   assign mem[434431:434400] = 32'b00000010111101001101110000001000;
   assign mem[434463:434432] = 32'b11110110011110110010011100000000;
   assign mem[434495:434464] = 32'b11100011111001000001000111000000;
   assign mem[434527:434496] = 32'b00000100100011000110110111000000;
   assign mem[434559:434528] = 32'b00000011100000000100011001011000;
   assign mem[434591:434560] = 32'b00000001100111100101110010100010;
   assign mem[434623:434592] = 32'b11111000011000010010011000111000;
   assign mem[434655:434624] = 32'b00000010111101000101110111101100;
   assign mem[434687:434656] = 32'b11111111010101111110111100110000;
   assign mem[434719:434688] = 32'b11110101111100001111000101000000;
   assign mem[434751:434720] = 32'b00000000101100111010110101101011;
   assign mem[434783:434752] = 32'b11111101101110100110100110111100;
   assign mem[434815:434784] = 32'b11110100101100001101101010000000;
   assign mem[434847:434816] = 32'b00000101010111001101101100100000;
   assign mem[434879:434848] = 32'b11111010010100001011001100111000;
   assign mem[434911:434880] = 32'b11111001010011010100110000101000;
   assign mem[434943:434912] = 32'b00000100100011101011110010010000;
   assign mem[434975:434944] = 32'b11111010011110100110000111111000;
   assign mem[435007:434976] = 32'b11111000011110111001100101000000;
   assign mem[435039:435008] = 32'b00000001101011101000001101100100;
   assign mem[435071:435040] = 32'b11111101111111000100100100101100;
   assign mem[435103:435072] = 32'b11111010101010010100010001001000;
   assign mem[435135:435104] = 32'b00000001110001101111101100101100;
   assign mem[435167:435136] = 32'b00000010111111110000010100101100;
   assign mem[435199:435168] = 32'b00000010010111010011100010010000;
   assign mem[435231:435200] = 32'b00000101110100101110110100001000;
   assign mem[435263:435232] = 32'b11111100101011000000001100010000;
   assign mem[435295:435264] = 32'b00000011110001010110011000101000;
   assign mem[435327:435296] = 32'b00000001011010111101110010110000;
   assign mem[435359:435328] = 32'b11111011001110001111101100001000;
   assign mem[435391:435360] = 32'b00000001101110000001110000000100;
   assign mem[435423:435392] = 32'b00000010110101101100011000011100;
   assign mem[435455:435424] = 32'b11110110000000100011110010010000;
   assign mem[435487:435456] = 32'b00000001111101111100100010100110;
   assign mem[435519:435488] = 32'b11111011101111110110111010011000;
   assign mem[435551:435520] = 32'b00000100100111000111010011000000;
   assign mem[435583:435552] = 32'b11111111000000101100000101100100;
   assign mem[435615:435584] = 32'b11111111011111101110111011111001;
   assign mem[435647:435616] = 32'b11111101101110010000101010100100;
   assign mem[435679:435648] = 32'b11110100010010110101101010100000;
   assign mem[435711:435680] = 32'b00000001100010001010001111111110;
   assign mem[435743:435712] = 32'b00000001101101011111011001010110;
   assign mem[435775:435744] = 32'b00000000101010010001100000011110;
   assign mem[435807:435776] = 32'b00000010111110010100000110110100;
   assign mem[435839:435808] = 32'b11110100010100010111110100010000;
   assign mem[435871:435840] = 32'b00000100110110100001111001110000;
   assign mem[435903:435872] = 32'b00000010110000001000110100110100;
   assign mem[435935:435904] = 32'b00000101010010001010111001110000;
   assign mem[435967:435936] = 32'b11111101001100101111101000011000;
   assign mem[435999:435968] = 32'b00000000100100000101010010010110;
   assign mem[436031:436000] = 32'b11111101110000001011100000010100;
   assign mem[436063:436032] = 32'b11111100001001111110010001101100;
   assign mem[436095:436064] = 32'b11111010111101010101001011011000;
   assign mem[436127:436096] = 32'b11111110000110110110011001000100;
   assign mem[436159:436128] = 32'b11111100001101101101110110110100;
   assign mem[436191:436160] = 32'b00000111100110010010001001101000;
   assign mem[436223:436192] = 32'b00000101011011001011011010111000;
   assign mem[436255:436224] = 32'b11111100001010001011001111100000;
   assign mem[436287:436256] = 32'b00000100110011010100000100011000;
   assign mem[436319:436288] = 32'b00000010001000010110011011111100;
   assign mem[436351:436320] = 32'b00000100100100111010000000011000;
   assign mem[436383:436352] = 32'b11100111010100111111010010000000;
   assign mem[436415:436384] = 32'b11111111000001000001110001010111;
   assign mem[436447:436416] = 32'b00000000001011101010100010101111;
   assign mem[436479:436448] = 32'b11111100001001001000100001001000;
   assign mem[436511:436480] = 32'b00000101001010100001100001011000;
   assign mem[436543:436512] = 32'b00000010101000110010110000100000;
   assign mem[436575:436544] = 32'b00000001001001000110000010110100;
   assign mem[436607:436576] = 32'b11101101111101010000110001000000;
   assign mem[436639:436608] = 32'b11111111000110010011100100110100;
   assign mem[436671:436640] = 32'b11110110010100011001101100100000;
   assign mem[436703:436672] = 32'b00000000110010011101111000011001;
   assign mem[436735:436704] = 32'b00000010101000010011000111111100;
   assign mem[436767:436736] = 32'b00000010100110110010000101111000;
   assign mem[436799:436768] = 32'b11110110001111011110101100110000;
   assign mem[436831:436800] = 32'b11111101011111101001101000011000;
   assign mem[436863:436832] = 32'b00000001111111010100011011101110;
   assign mem[436895:436864] = 32'b11111011001001100110000011011000;
   assign mem[436927:436896] = 32'b00001000001001111011011011100000;
   assign mem[436959:436928] = 32'b11111010100110101110000100011000;
   assign mem[436991:436960] = 32'b00000101100101010110100111010000;
   assign mem[437023:436992] = 32'b11110110010011011011100100010000;
   assign mem[437055:437024] = 32'b11111000100010001111101110101000;
   assign mem[437087:437056] = 32'b11111011011011101111001101001000;
   assign mem[437119:437088] = 32'b00000000001010010010101011100000;
   assign mem[437151:437120] = 32'b11111010100101110100111100100000;
   assign mem[437183:437152] = 32'b00000100101000101001011100111000;
   assign mem[437215:437184] = 32'b11111000011100000101010111100000;
   assign mem[437247:437216] = 32'b11110110100001110011001101010000;
   assign mem[437279:437248] = 32'b00001001001001000111101011110000;
   assign mem[437311:437280] = 32'b00000111000010011111111101101000;
   assign mem[437343:437312] = 32'b11110110010000111101011010100000;
   assign mem[437375:437344] = 32'b00000110001001111010100000101000;
   assign mem[437407:437376] = 32'b11111000110100101001011101001000;
   assign mem[437439:437408] = 32'b00000111001110100011110111110000;
   assign mem[437471:437440] = 32'b00000010000111001110001001111000;
   assign mem[437503:437472] = 32'b11111010000101110010000001001000;
   assign mem[437535:437504] = 32'b00000001111010111110000011011110;
   assign mem[437567:437536] = 32'b11111111110000111110001111101100;
   assign mem[437599:437568] = 32'b11110110010011011010011100010000;
   assign mem[437631:437600] = 32'b11111110110001010100110111011010;
   assign mem[437663:437632] = 32'b00000010001010010111101011011100;
   assign mem[437695:437664] = 32'b11110011100001000110000100110000;
   assign mem[437727:437696] = 32'b00000011000011110100100101100000;
   assign mem[437759:437728] = 32'b11110110000111111010101011010000;
   assign mem[437791:437760] = 32'b00000010011000011111100011001100;
   assign mem[437823:437792] = 32'b11110001001110100100011100010000;
   assign mem[437855:437824] = 32'b00000100100000110011101100011000;
   assign mem[437887:437856] = 32'b11111111111111000001000011011010;
   assign mem[437919:437888] = 32'b11110101001110110001001001000000;
   assign mem[437951:437920] = 32'b00000011110111000101000101111000;
   assign mem[437983:437952] = 32'b00000010000101100000001010101100;
   assign mem[438015:437984] = 32'b11110000001010100010001100000000;
   assign mem[438047:438016] = 32'b00000110011001010110111101010000;
   assign mem[438079:438048] = 32'b11111000110011101101111111001000;
   assign mem[438111:438080] = 32'b11111101111010001011001101000000;
   assign mem[438143:438112] = 32'b00010111000101101101001001100000;
   assign mem[438175:438144] = 32'b00000011010011111010010000101000;
   assign mem[438207:438176] = 32'b11111000011011111100111011010000;
   assign mem[438239:438208] = 32'b00000001011100001001100100001110;
   assign mem[438271:438240] = 32'b00001001101111101001001011110000;
   assign mem[438303:438272] = 32'b11110011000000000110111001000000;
   assign mem[438335:438304] = 32'b00001010110010100110100000110000;
   assign mem[438367:438336] = 32'b11111110001001010100010100011000;
   assign mem[438399:438368] = 32'b11110010110101100100101000100000;
   assign mem[438431:438400] = 32'b00001011000001110011101101010000;
   assign mem[438463:438432] = 32'b11111101100010101100101111101000;
   assign mem[438495:438464] = 32'b00000000110100100001001011101111;
   assign mem[438527:438496] = 32'b11111010011001110101011101011000;
   assign mem[438559:438528] = 32'b11111011110100100010010001010000;
   assign mem[438591:438560] = 32'b11111111110101110010011001100110;
   assign mem[438623:438592] = 32'b00000100010011110111110000011000;
   assign mem[438655:438624] = 32'b11111011101010100110111000010000;
   assign mem[438687:438656] = 32'b00001000111110011000001110000000;
   assign mem[438719:438688] = 32'b11101011110100011010010101000000;
   assign mem[438751:438720] = 32'b11100110011111000000011011100000;
   assign mem[438783:438752] = 32'b00000100010100111001110111100000;
   assign mem[438815:438784] = 32'b00000011001111000110111111110100;
   assign mem[438847:438816] = 32'b00000110111111111001000100001000;
   assign mem[438879:438848] = 32'b11111110010111001000101101110110;
   assign mem[438911:438880] = 32'b00001001111101111111001011010000;
   assign mem[438943:438912] = 32'b11101100100110111111100111100000;
   assign mem[438975:438944] = 32'b00000000001101100111010101011000;
   assign mem[439007:438976] = 32'b11111001100011011000110110100000;
   assign mem[439039:439008] = 32'b00000100000111111011101010010000;
   assign mem[439071:439040] = 32'b00000001101000111001010001111100;
   assign mem[439103:439072] = 32'b00000101000111010011011000100000;
   assign mem[439135:439104] = 32'b00000000010011111110110010100011;
   assign mem[439167:439136] = 32'b11111101011110011111100001000000;
   assign mem[439199:439168] = 32'b11111010110010101101110111100000;
   assign mem[439231:439200] = 32'b11111100110100100101101100010100;
   assign mem[439263:439232] = 32'b00000001011111101010110000000110;
   assign mem[439295:439264] = 32'b11110111010110100011101011000000;
   assign mem[439327:439296] = 32'b00000010010101101000010001110100;
   assign mem[439359:439328] = 32'b00000001111111101101111000000100;
   assign mem[439391:439360] = 32'b11111010101110000100110100100000;
   assign mem[439423:439392] = 32'b00001101100101100000110001010000;
   assign mem[439455:439424] = 32'b11110011110000100010011011110000;
   assign mem[439487:439456] = 32'b00001000100001111101000011100000;
   assign mem[439519:439488] = 32'b11110000111010000111111001010000;
   assign mem[439551:439520] = 32'b00001011100100011010010000010000;
   assign mem[439583:439552] = 32'b11101111010000011100100000000000;
   assign mem[439615:439584] = 32'b11110111100100000001010100000000;
   assign mem[439647:439616] = 32'b11101111010011001011101001100000;
   assign mem[439679:439648] = 32'b00000110101100101010001110111000;
   assign mem[439711:439680] = 32'b00000011111101100101001001001000;
   assign mem[439743:439712] = 32'b00010110000000001101010101000000;
   assign mem[439775:439744] = 32'b11111001000100111110100000000000;
   assign mem[439807:439776] = 32'b11110011101110110011011011100000;
   assign mem[439839:439808] = 32'b00000100101111000111000100101000;
   assign mem[439871:439840] = 32'b11111001110000101000100001010000;
   assign mem[439903:439872] = 32'b00000000011010000111001110101111;
   assign mem[439935:439904] = 32'b00000011100001101101110101011100;
   assign mem[439967:439936] = 32'b00000001010111010001111111111110;
   assign mem[439999:439968] = 32'b11111011100011111110000100011000;
   assign mem[440031:440000] = 32'b11111110100100001111100111101110;
   assign mem[440063:440032] = 32'b11111111010010011101101011011011;
   assign mem[440095:440064] = 32'b00000000001100110101001101101101;
   assign mem[440127:440096] = 32'b00000001100100001101010010111000;
   assign mem[440159:440128] = 32'b11111110010010111010100101010000;
   assign mem[440191:440160] = 32'b00000010001010101011110001111100;
   assign mem[440223:440192] = 32'b00000000111000101000100111110000;
   assign mem[440255:440224] = 32'b11111000100101111010110111010000;
   assign mem[440287:440256] = 32'b11111111011011001111001110101100;
   assign mem[440319:440288] = 32'b00000000101001010100110101100101;
   assign mem[440351:440320] = 32'b11111100001011101111111011000000;
   assign mem[440383:440352] = 32'b11111111011011001111000000110011;
   assign mem[440415:440384] = 32'b00000010101101000001110010111100;
   assign mem[440447:440416] = 32'b11111011101011010011100001010000;
   assign mem[440479:440448] = 32'b00000111001101101001011101011000;
   assign mem[440511:440480] = 32'b00000010010011000100100011100000;
   assign mem[440543:440512] = 32'b11110110101010010100001011100000;
   assign mem[440575:440544] = 32'b00000101001110011100100010111000;
   assign mem[440607:440576] = 32'b00000100110101010001110101111000;
   assign mem[440639:440608] = 32'b00000110010001010010001010010000;
   assign mem[440671:440640] = 32'b11111000101110010011001011110000;
   assign mem[440703:440672] = 32'b00000111000111011000101110101000;
   assign mem[440735:440704] = 32'b11111011110000011000111110010000;
   assign mem[440767:440736] = 32'b11110101010100000110100011110000;
   assign mem[440799:440768] = 32'b00001000111011001010110100100000;
   assign mem[440831:440800] = 32'b11110011100100111000101101100000;
   assign mem[440863:440832] = 32'b11111010110000000001011110010000;
   assign mem[440895:440864] = 32'b00000101101000110000010101011000;
   assign mem[440927:440896] = 32'b11111100101100101001110101101000;
   assign mem[440959:440928] = 32'b00000100011100001111110011010000;
   assign mem[440991:440960] = 32'b00000010011100011101000011100000;
   assign mem[441023:440992] = 32'b00000001011101100110100011110010;
   assign mem[441055:441024] = 32'b11111110010001101010100010101110;
   assign mem[441087:441056] = 32'b11111110001001100101001111100000;
   assign mem[441119:441088] = 32'b11111111101000011101101101111000;
   assign mem[441151:441120] = 32'b00000000011111010011011100000000;
   assign mem[441183:441152] = 32'b00000000010111100110001000001100;
   assign mem[441215:441184] = 32'b11111001111011111010001111110000;
   assign mem[441247:441216] = 32'b11111110000100000011000101101110;
   assign mem[441279:441248] = 32'b11111111101001101010110110001000;
   assign mem[441311:441280] = 32'b11101100011011010110111100000000;
   assign mem[441343:441312] = 32'b00001101110110100010011101000000;
   assign mem[441375:441344] = 32'b00000110011011010101110110001000;
   assign mem[441407:441376] = 32'b00001010011010110110100010100000;
   assign mem[441439:441408] = 32'b11111011011100111101101010101000;
   assign mem[441471:441440] = 32'b00000111010011010011000100011000;
   assign mem[441503:441472] = 32'b11101110000111100000011001100000;
   assign mem[441535:441504] = 32'b00001001010111011001110110010000;
   assign mem[441567:441536] = 32'b11101101110010011010101100100000;
   assign mem[441599:441568] = 32'b11111010110110111110011000010000;
   assign mem[441631:441600] = 32'b11111111000010001010011010001010;
   assign mem[441663:441632] = 32'b11111010011100000010110010000000;
   assign mem[441695:441664] = 32'b00000000101000011000011110101010;
   assign mem[441727:441696] = 32'b11111100101001000101101100001100;
   assign mem[441759:441728] = 32'b11111001100110111010111111001000;
   assign mem[441791:441760] = 32'b00000010110100111011001100111100;
   assign mem[441823:441792] = 32'b11111001100001001111001011110000;
   assign mem[441855:441824] = 32'b11111001011001000111100110001000;
   assign mem[441887:441856] = 32'b11111101101100110101001100100100;
   assign mem[441919:441888] = 32'b11111111101010100100010111100111;
   assign mem[441951:441920] = 32'b00000011100001101110100010111000;
   assign mem[441983:441952] = 32'b00001001110010001110010011010000;
   assign mem[442015:441984] = 32'b11111110111000100100011010110110;
   assign mem[442047:442016] = 32'b00000011000110011000010000110000;
   assign mem[442079:442048] = 32'b11111010011111110100010011111000;
   assign mem[442111:442080] = 32'b00000101110111111000101101100000;
   assign mem[442143:442112] = 32'b11110010101000110001011000000000;
   assign mem[442175:442144] = 32'b11110000111000001100111001100000;
   assign mem[442207:442176] = 32'b11111100010100110101101100111100;
   assign mem[442239:442208] = 32'b00000010000101010111011011010000;
   assign mem[442271:442240] = 32'b00000010001100010110111010011000;
   assign mem[442303:442272] = 32'b11111100001001000001101000110100;
   assign mem[442335:442304] = 32'b00000000010011100000110101000101;
   assign mem[442367:442336] = 32'b11111111101101100011100100110100;
   assign mem[442399:442368] = 32'b11110111101110111001111011110000;
   assign mem[442431:442400] = 32'b11111111110000000111111100010100;
   assign mem[442463:442432] = 32'b11111110110001011001010000001100;
   assign mem[442495:442464] = 32'b11111000001111010110110010101000;
   assign mem[442527:442496] = 32'b00000010110011100011010101000100;
   assign mem[442559:442528] = 32'b00000100000100000100001111100000;
   assign mem[442591:442560] = 32'b11110101100101110000110010010000;
   assign mem[442623:442592] = 32'b11111100001000100101000001100100;
   assign mem[442655:442624] = 32'b00000010001000111111110010100100;
   assign mem[442687:442656] = 32'b00000100100110000101000101011000;
   assign mem[442719:442688] = 32'b11111111010011110010001101101101;
   assign mem[442751:442720] = 32'b00001010110011100100000111100000;
   assign mem[442783:442752] = 32'b11110101011011100110010111000000;
   assign mem[442815:442784] = 32'b11111111011000011101001001111010;
   assign mem[442847:442816] = 32'b11110001110111000101101011100000;
   assign mem[442879:442848] = 32'b00000011000010000100100100010100;
   assign mem[442911:442880] = 32'b00000101010010110000101101011000;
   assign mem[442943:442912] = 32'b11110110010111001101101011100000;
   assign mem[442975:442944] = 32'b00000011000100110011111100110000;
   assign mem[443007:442976] = 32'b11111110111001000101000000001110;
   assign mem[443039:443008] = 32'b11111000100101001000100001110000;
   assign mem[443071:443040] = 32'b11111111101011001010000110010100;
   assign mem[443103:443072] = 32'b00000101101110110100100011001000;
   assign mem[443135:443104] = 32'b11111101011110100110010101010100;
   assign mem[443167:443136] = 32'b00000001100101100001001111110010;
   assign mem[443199:443168] = 32'b11111111001000100100101110000011;
   assign mem[443231:443200] = 32'b00000000001111011011011110100110;
   assign mem[443263:443232] = 32'b11111101111100110100110011000000;
   assign mem[443295:443264] = 32'b00000011001011111111101011000100;
   assign mem[443327:443296] = 32'b11111111100100001101111001111111;
   assign mem[443359:443328] = 32'b11111011110101100100000001011000;
   assign mem[443391:443360] = 32'b00000001001011111001001001001100;
   assign mem[443423:443392] = 32'b00000000101101100011000101000111;
   assign mem[443455:443424] = 32'b11111011000110100110111010001000;
   assign mem[443487:443456] = 32'b11111010001000111110000010100000;
   assign mem[443519:443488] = 32'b00000001001101001011011111000100;
   assign mem[443551:443520] = 32'b11111111010011100111011011010101;
   assign mem[443583:443552] = 32'b11111011110111001100010110101000;
   assign mem[443615:443584] = 32'b11111110010110101100111000010000;
   assign mem[443647:443616] = 32'b11111110101101000101111011110010;
   assign mem[443679:443648] = 32'b11111101011011011001001101001100;
   assign mem[443711:443680] = 32'b00000010000101111001101001111100;
   assign mem[443743:443712] = 32'b00000010110110000001011111000000;
   assign mem[443775:443744] = 32'b11111101110011111011110010010000;
   assign mem[443807:443776] = 32'b11111100111101001010011011100000;
   assign mem[443839:443808] = 32'b00000010101011100000000110000100;
   assign mem[443871:443840] = 32'b00001001111011001101111101110000;
   assign mem[443903:443872] = 32'b11111010100110100000010011110000;
   assign mem[443935:443904] = 32'b00000111101001100110111101010000;
   assign mem[443967:443936] = 32'b00000000011010111010110000100011;
   assign mem[443999:443968] = 32'b11110111110010011111000110110000;
   assign mem[444031:444000] = 32'b00000011001011111011000001010100;
   assign mem[444063:444032] = 32'b11111111001010001011011111011000;
   assign mem[444095:444064] = 32'b11110101010011000001101111010000;
   assign mem[444127:444096] = 32'b11111001000011100010111111100000;
   assign mem[444159:444128] = 32'b11111011011000011110111010011000;
   assign mem[444191:444160] = 32'b00000010111101111100000100110100;
   assign mem[444223:444192] = 32'b11111011111101110011100000110000;
   assign mem[444255:444224] = 32'b00000100000001101111001110101000;
   assign mem[444287:444256] = 32'b11111111110001111100000100010111;
   assign mem[444319:444288] = 32'b11111001110111011110111111100000;
   assign mem[444351:444320] = 32'b11111101010010011101100011010000;
   assign mem[444383:444352] = 32'b00000011000110010111101010011000;
   assign mem[444415:444384] = 32'b11101110010010000010011110000000;
   assign mem[444447:444416] = 32'b00000101010000000101111000011000;
   assign mem[444479:444448] = 32'b11111100011111100110010100101100;
   assign mem[444511:444480] = 32'b00001011001000110011101100000000;
   assign mem[444543:444512] = 32'b11110011010111111110101001010000;
   assign mem[444575:444544] = 32'b11111111011000101010101100101111;
   assign mem[444607:444576] = 32'b00000011100010110101010111011100;
   assign mem[444639:444608] = 32'b00000100001001100011001101010000;
   assign mem[444671:444640] = 32'b00000101100001001011100000011000;
   assign mem[444703:444672] = 32'b11111010110001000100001100011000;
   assign mem[444735:444704] = 32'b00000011000101001110110110111100;
   assign mem[444767:444736] = 32'b11111101011000001001110001001000;
   assign mem[444799:444768] = 32'b11111001100110000110001001111000;
   assign mem[444831:444800] = 32'b00000101010001011000011100010000;
   assign mem[444863:444832] = 32'b00000101011111100001010000000000;
   assign mem[444895:444864] = 32'b11111011001011110101011101010000;
   assign mem[444927:444896] = 32'b11110101010001110000110110100000;
   assign mem[444959:444928] = 32'b11111110101010000101110111101000;
   assign mem[444991:444960] = 32'b11111011010111100110000000110000;
   assign mem[445023:444992] = 32'b00000101111111000100011100111000;
   assign mem[445055:445024] = 32'b00000100010111100011000101010000;
   assign mem[445087:445056] = 32'b00000010011010111000101110101000;
   assign mem[445119:445088] = 32'b11111011110100111101001011100000;
   assign mem[445151:445120] = 32'b00000010111110011001001000000100;
   assign mem[445183:445152] = 32'b11111110010001101011010011010000;
   assign mem[445215:445184] = 32'b00000010111110110000010100100000;
   assign mem[445247:445216] = 32'b11111110101111001100001100101110;
   assign mem[445279:445248] = 32'b11111101000011100101101110101100;
   assign mem[445311:445280] = 32'b00000011011110000110010001001000;
   assign mem[445343:445312] = 32'b00000001010000100001100110110010;
   assign mem[445375:445344] = 32'b00000001011100010100000100011000;
   assign mem[445407:445376] = 32'b00000000100111001001011111001110;
   assign mem[445439:445408] = 32'b11111101100000111011110000010000;
   assign mem[445471:445440] = 32'b00001000000000011001100010000000;
   assign mem[445503:445472] = 32'b11111011101001001110010101110000;
   assign mem[445535:445504] = 32'b00000101110010001001000000011000;
   assign mem[445567:445536] = 32'b11111111100100000000110000000100;
   assign mem[445599:445568] = 32'b00000010111010011000001011110000;
   assign mem[445631:445600] = 32'b00000010110111110010001111011000;
   assign mem[445663:445632] = 32'b11111110110101010011110100111000;
   assign mem[445695:445664] = 32'b11110111111111111100110111100000;
   assign mem[445727:445696] = 32'b11111001011000010111100111111000;
   assign mem[445759:445728] = 32'b11111001111101111001100001100000;
   assign mem[445791:445760] = 32'b11110001111110101010110011010000;
   assign mem[445823:445792] = 32'b11111110001011000101000110000000;
   assign mem[445855:445824] = 32'b00000010000100111110111110111000;
   assign mem[445887:445856] = 32'b11111110110101100100100100000100;
   assign mem[445919:445888] = 32'b11111101101000001101001110000000;
   assign mem[445951:445920] = 32'b00000000100101001000011110010111;
   assign mem[445983:445952] = 32'b11111001100100011011111011110000;
   assign mem[446015:445984] = 32'b11111111011101101101110011110011;
   assign mem[446047:446016] = 32'b11111100011000111000110111100100;
   assign mem[446079:446048] = 32'b00000101110001001111000001010000;
   assign mem[446111:446080] = 32'b00000101001010101010100011010000;
   assign mem[446143:446112] = 32'b11111111000101001010001100001100;
   assign mem[446175:446144] = 32'b11111101110000111111001011111000;
   assign mem[446207:446176] = 32'b11111100000001111110101110100000;
   assign mem[446239:446208] = 32'b00000110011111100001110011100000;
   assign mem[446271:446240] = 32'b11111011100101010100010110011000;
   assign mem[446303:446272] = 32'b11111100100011010000011010101000;
   assign mem[446335:446304] = 32'b00000101100100010000000111001000;
   assign mem[446367:446336] = 32'b11111100100101100000110000000000;
   assign mem[446399:446368] = 32'b00000011101010110000000111110000;
   assign mem[446431:446400] = 32'b00000011101000101101000111100000;
   assign mem[446463:446432] = 32'b00000100100101011101100111011000;
   assign mem[446495:446464] = 32'b00000011110000101000101001100100;
   assign mem[446527:446496] = 32'b11111111101010000110010000011011;
   assign mem[446559:446528] = 32'b00000010000000101010001001001000;
   assign mem[446591:446560] = 32'b11111110100011011011001000000010;
   assign mem[446623:446592] = 32'b00000010010100111001111000100100;
   assign mem[446655:446624] = 32'b11111010101011100101011101000000;
   assign mem[446687:446656] = 32'b00000010110000100001010101110100;
   assign mem[446719:446688] = 32'b11111010110011101100000100101000;
   assign mem[446751:446720] = 32'b00000100110000110111001011010000;
   assign mem[446783:446752] = 32'b00000011100011101111001010110100;
   assign mem[446815:446784] = 32'b00000011011001010110101110000100;
   assign mem[446847:446816] = 32'b00000001101110000110010101111000;
   assign mem[446879:446848] = 32'b11111110011100000010010101110010;
   assign mem[446911:446880] = 32'b00000011100100101100001100000000;
   assign mem[446943:446912] = 32'b00000010111111111100010011010100;
   assign mem[446975:446944] = 32'b11110100101111011110000100110000;
   assign mem[447007:446976] = 32'b00000010110000101001011110010000;
   assign mem[447039:447008] = 32'b11111010111111100100000110001000;
   assign mem[447071:447040] = 32'b11111111010101001100100011111110;
   assign mem[447103:447072] = 32'b00000101110000110111110000011000;
   assign mem[447135:447104] = 32'b00000000001111010011100111100101;
   assign mem[447167:447136] = 32'b11111111011100101110001001111000;
   assign mem[447199:447168] = 32'b11111011100000001111111000100000;
   assign mem[447231:447200] = 32'b00000011100011111000000011011100;
   assign mem[447263:447232] = 32'b11111100101100000001010001111100;
   assign mem[447295:447264] = 32'b11111110111010111111100001001110;
   assign mem[447327:447296] = 32'b00000010101111011100011111000000;
   assign mem[447359:447328] = 32'b11111110000001010100101101100000;
   assign mem[447391:447360] = 32'b11111111111111111010001100101010;
   assign mem[447423:447392] = 32'b00000000101111111101100111001111;
   assign mem[447455:447424] = 32'b00000110110111000010000111111000;
   assign mem[447487:447456] = 32'b11111110001011001101000000111010;
   assign mem[447519:447488] = 32'b11111010011011010000010011000000;
   assign mem[447551:447520] = 32'b00000100110001000000110100001000;
   assign mem[447583:447552] = 32'b11111111010011110011111110111100;
   assign mem[447615:447584] = 32'b11110110110100110101101101000000;
   assign mem[447647:447616] = 32'b11111110110001100111010111101110;
   assign mem[447679:447648] = 32'b11111101001110110110101111101100;
   assign mem[447711:447680] = 32'b00000100011000100110010110001000;
   assign mem[447743:447712] = 32'b00001101010011100011011011100000;
   assign mem[447775:447744] = 32'b11111100010100111011110110001000;
   assign mem[447807:447776] = 32'b11110101110000001010000110110000;
   assign mem[447839:447808] = 32'b00000010100110111110011001000000;
   assign mem[447871:447840] = 32'b11111000100000111000101100110000;
   assign mem[447903:447872] = 32'b11110110101100001111111011000000;
   assign mem[447935:447904] = 32'b00000110111110110001010110000000;
   assign mem[447967:447936] = 32'b11111110111111111000010001101000;
   assign mem[447999:447968] = 32'b00000110011110101000100001011000;
   assign mem[448031:448000] = 32'b00000100000110001011010111111000;
   assign mem[448063:448032] = 32'b00000000110011110100100010000101;
   assign mem[448095:448064] = 32'b00000011011010110111110111010000;
   assign mem[448127:448096] = 32'b00000100000011100110010100110000;
   assign mem[448159:448128] = 32'b11111001001000011011110001101000;
   assign mem[448191:448160] = 32'b00000100010000110001001010010000;
   assign mem[448223:448192] = 32'b11111111101110101011100101001100;
   assign mem[448255:448224] = 32'b00000101001001111001100011010000;
   assign mem[448287:448256] = 32'b00000010010100110000010111111000;
   assign mem[448319:448288] = 32'b11111001011101111110001011010000;
   assign mem[448351:448320] = 32'b00000001110100110001101000001000;
   assign mem[448383:448352] = 32'b11111011101100100100110010110000;
   assign mem[448415:448384] = 32'b11111101111001011100100001100100;
   assign mem[448447:448416] = 32'b00000000101111100011001110010001;
   assign mem[448479:448448] = 32'b11111100100001010001101110101100;
   assign mem[448511:448480] = 32'b00000010000111100101001101001100;
   assign mem[448543:448512] = 32'b00000011001111000110001011111100;
   assign mem[448575:448544] = 32'b11111110100110011111110011100110;
   assign mem[448607:448576] = 32'b11111110011111010011011100110000;
   assign mem[448639:448608] = 32'b00000000101100010010110101100101;
   assign mem[448671:448640] = 32'b00000000000010010101010011010110;
   assign mem[448703:448672] = 32'b00000101010100110000000111000000;
   assign mem[448735:448704] = 32'b11110111001101011110100100000000;
   assign mem[448767:448736] = 32'b00001010011111010111100011100000;
   assign mem[448799:448768] = 32'b11110010101110101100111110010000;
   assign mem[448831:448800] = 32'b00001000110011001010001100000000;
   assign mem[448863:448832] = 32'b11111000100101111100010001101000;
   assign mem[448895:448864] = 32'b11101111001010011010111101000000;
   assign mem[448927:448896] = 32'b11110001010101010000101101100000;
   assign mem[448959:448928] = 32'b00001000001010011111111101010000;
   assign mem[448991:448960] = 32'b00001001001011000010101011010000;
   assign mem[449023:448992] = 32'b11111001110000001001111000110000;
   assign mem[449055:449024] = 32'b00000101001011100001100101101000;
   assign mem[449087:449056] = 32'b00000010101100000111010000001100;
   assign mem[449119:449088] = 32'b11111000110100011101000100010000;
   assign mem[449151:449120] = 32'b00000100110100001010011111000000;
   assign mem[449183:449152] = 32'b11111110101010010010011010010010;
   assign mem[449215:449184] = 32'b11110100111010110111001100100000;
   assign mem[449247:449216] = 32'b11110011110010110110011001010000;
   assign mem[449279:449248] = 32'b00000010101110010110010011100000;
   assign mem[449311:449280] = 32'b11101000001110111010001111100000;
   assign mem[449343:449312] = 32'b00000100100101001100010101000000;
   assign mem[449375:449344] = 32'b11111110000101010001010110001110;
   assign mem[449407:449376] = 32'b00001010110001101111010110000000;
   assign mem[449439:449408] = 32'b00000010110010001001011111111100;
   assign mem[449471:449440] = 32'b00001111001110100100100110010000;
   assign mem[449503:449472] = 32'b11101101100110111110100000100000;
   assign mem[449535:449504] = 32'b11111111110110101101010100110110;
   assign mem[449567:449536] = 32'b11101010100111010001100001100000;
   assign mem[449599:449568] = 32'b00000101101001101011110011101000;
   assign mem[449631:449600] = 32'b11110011011111111010001101000000;
   assign mem[449663:449632] = 32'b00000001010011010111010000001000;
   assign mem[449695:449664] = 32'b11111110000111010010000111000110;
   assign mem[449727:449696] = 32'b11111000011110110110101101000000;
   assign mem[449759:449728] = 32'b00000101001100111001101011110000;
   assign mem[449791:449760] = 32'b11111111100101100001100101100001;
   assign mem[449823:449792] = 32'b11111000100000010011110011101000;
   assign mem[449855:449824] = 32'b00000111101111001100000001111000;
   assign mem[449887:449856] = 32'b11111010110111110101000000000000;
   assign mem[449919:449888] = 32'b00000110000001001100101011101000;
   assign mem[449951:449920] = 32'b00001000101011000111010110000000;
   assign mem[449983:449952] = 32'b00000010000001101011101000111000;
   assign mem[450015:449984] = 32'b00000101111011000000000011111000;
   assign mem[450047:450016] = 32'b11111111100101100001101111011111;
   assign mem[450079:450048] = 32'b11111011011111000101001010100000;
   assign mem[450111:450080] = 32'b11111110110101101110010011111000;
   assign mem[450143:450112] = 32'b11111110111000100001111011011000;
   assign mem[450175:450144] = 32'b11111101101011000011001001001000;
   assign mem[450207:450176] = 32'b00000110100101001011110111101000;
   assign mem[450239:450208] = 32'b11111011011011110001010000000000;
   assign mem[450271:450240] = 32'b00000011100010110111001101000000;
   assign mem[450303:450272] = 32'b00000101011000011110100011001000;
   assign mem[450335:450304] = 32'b11111111110110000000111000011010;
   assign mem[450367:450336] = 32'b11101111011010100111011111100000;
   assign mem[450399:450368] = 32'b11111110000101101011100110110010;
   assign mem[450431:450400] = 32'b11110100001011010011110111010000;
   assign mem[450463:450432] = 32'b11111001110011111010010000101000;
   assign mem[450495:450464] = 32'b00000000101100100001011011111101;
   assign mem[450527:450496] = 32'b00000100000011111110011101111000;
   assign mem[450559:450528] = 32'b00000000001110010001000010110111;
   assign mem[450591:450560] = 32'b00000110011101011001100110101000;
   assign mem[450623:450592] = 32'b11110101111101111001011111000000;
   assign mem[450655:450624] = 32'b11111011101010010010100001000000;
   assign mem[450687:450656] = 32'b11111010110111001100010001100000;
   assign mem[450719:450688] = 32'b11111110011100001000000100010000;
   assign mem[450751:450720] = 32'b11111011100011011001100100001000;
   assign mem[450783:450752] = 32'b11111110000000011001111001000100;
   assign mem[450815:450784] = 32'b11111111101000111111111010001000;
   assign mem[450847:450816] = 32'b00000010100010111110000111010000;
   assign mem[450879:450848] = 32'b00000110011101010101101100110000;
   assign mem[450911:450880] = 32'b00001111101000101010110111110000;
   assign mem[450943:450912] = 32'b00001100111010001010011010000000;
   assign mem[450975:450944] = 32'b11100010001010110101110100000000;
   assign mem[451007:450976] = 32'b00000001000110100011001010101100;
   assign mem[451039:451008] = 32'b11111011001000001111001100010000;
   assign mem[451071:451040] = 32'b00000010110100111110011101001000;
   assign mem[451103:451072] = 32'b00000000010011011110001101001111;
   assign mem[451135:451104] = 32'b00000100011110101011110001011000;
   assign mem[451167:451136] = 32'b11110011001011111110001010110000;
   assign mem[451199:451168] = 32'b00000100010010100011000101001000;
   assign mem[451231:451200] = 32'b00000111000011000111011111000000;
   assign mem[451263:451232] = 32'b11111010011000111000011010000000;
   assign mem[451295:451264] = 32'b00000110110110010011000011110000;
   assign mem[451327:451296] = 32'b00000100010011001101100011001000;
   assign mem[451359:451328] = 32'b11110100010011101111101110100000;
   assign mem[451391:451360] = 32'b00000001000011101001101101011010;
   assign mem[451423:451392] = 32'b00000111000110001010000110010000;
   assign mem[451455:451424] = 32'b11110100010010000110110011000000;
   assign mem[451487:451456] = 32'b00000011101001111110011110111000;
   assign mem[451519:451488] = 32'b11111110110010001000101011111100;
   assign mem[451551:451520] = 32'b11111101110100001100001101101000;
   assign mem[451583:451552] = 32'b11111110010010111000011100000110;
   assign mem[451615:451584] = 32'b11111100100010110000101011110100;
   assign mem[451647:451616] = 32'b00000000101111111001110010000111;
   assign mem[451679:451648] = 32'b11111101010010010110011000111000;
   assign mem[451711:451680] = 32'b11111111111000110111101001110100;
   assign mem[451743:451712] = 32'b00000011000010100110111000011100;
   assign mem[451775:451744] = 32'b11111010011111100010110001011000;
   assign mem[451807:451776] = 32'b11111111101111011101011110111110;
   assign mem[451839:451808] = 32'b11111110001111010111010110100100;
   assign mem[451871:451840] = 32'b00000000101110001111100111000001;
   assign mem[451903:451872] = 32'b11111010110111111100000100100000;
   assign mem[451935:451904] = 32'b00000111010111011101010011100000;
   assign mem[451967:451936] = 32'b00000000011111100011000101010010;
   assign mem[451999:451968] = 32'b11111011001111111000110110000000;
   assign mem[452031:452000] = 32'b00000010100101111110100011000100;
   assign mem[452063:452032] = 32'b00000011000010100100110001011000;
   assign mem[452095:452064] = 32'b11110111010100010110011000100000;
   assign mem[452127:452096] = 32'b11110111100110100000000111010000;
   assign mem[452159:452128] = 32'b11111111101001110001101101110110;
   assign mem[452191:452160] = 32'b00000010110000010010000111011000;
   assign mem[452223:452192] = 32'b00000000111101010010110100101111;
   assign mem[452255:452224] = 32'b11111011000101001100100100010000;
   assign mem[452287:452256] = 32'b00000000001000100110011011101001;
   assign mem[452319:452288] = 32'b00000100111110111000010110111000;
   assign mem[452351:452320] = 32'b11111110001011010111001010000000;
   assign mem[452383:452352] = 32'b11111101101101001110101111010000;
   assign mem[452415:452384] = 32'b00000101000010101110000010100000;
   assign mem[452447:452416] = 32'b11110111101010011010001100010000;
   assign mem[452479:452448] = 32'b00000010101100111011100100111000;
   assign mem[452511:452480] = 32'b11111000010011010101100001101000;
   assign mem[452543:452512] = 32'b00001010001100111010101110000000;
   assign mem[452575:452544] = 32'b11111100011110011100010010110000;
   assign mem[452607:452576] = 32'b11110001011011000000111101110000;
   assign mem[452639:452608] = 32'b00000100111110110001010000010000;
   assign mem[452671:452640] = 32'b00000111101011111110011011010000;
   assign mem[452703:452672] = 32'b11110011011101000111101010100000;
   assign mem[452735:452704] = 32'b00000100010111111111111101101000;
   assign mem[452767:452736] = 32'b11111101000001110110001010010000;
   assign mem[452799:452768] = 32'b00001001101011101011110101110000;
   assign mem[452831:452800] = 32'b00000111100110110000011111100000;
   assign mem[452863:452832] = 32'b11111100010111110110011001000000;
   assign mem[452895:452864] = 32'b11111110010010101001100101010100;
   assign mem[452927:452896] = 32'b00000011000011001011111010100100;
   assign mem[452959:452928] = 32'b00000001110000110110010110010110;
   assign mem[452991:452960] = 32'b00000100101110001011100100111000;
   assign mem[453023:452992] = 32'b11111110110010000000100000111110;
   assign mem[453055:453024] = 32'b11111110100011011000110110101100;
   assign mem[453087:453056] = 32'b11111001000111100001111101010000;
   assign mem[453119:453088] = 32'b00000010000100111001101010111000;
   assign mem[453151:453120] = 32'b11111110111101100010111000100100;
   assign mem[453183:453152] = 32'b00001101110100011111100111010000;
   assign mem[453215:453184] = 32'b11101110000000101100100000100000;
   assign mem[453247:453216] = 32'b11111111011101111010111001101111;
   assign mem[453279:453248] = 32'b11100110111101001001111101100000;
   assign mem[453311:453280] = 32'b00000100001010000100001011101000;
   assign mem[453343:453312] = 32'b00000011011011110111011110001100;
   assign mem[453375:453344] = 32'b11110111110000011101001011100000;
   assign mem[453407:453376] = 32'b11110111111010011101110101010000;
   assign mem[453439:453408] = 32'b00000101000000111000010100001000;
   assign mem[453471:453440] = 32'b11100110000110100110100110100000;
   assign mem[453503:453472] = 32'b00000101011100001100101001001000;
   assign mem[453535:453504] = 32'b00000000001011000101111010101001;
   assign mem[453567:453536] = 32'b11110111000110100100001100000000;
   assign mem[453599:453568] = 32'b00000011001110011000110001101000;
   assign mem[453631:453600] = 32'b11111001101011011000100111100000;
   assign mem[453663:453632] = 32'b11100100111000101011000010000000;
   assign mem[453695:453664] = 32'b00000110010110110011010000111000;
   assign mem[453727:453696] = 32'b11111010011001001010100101110000;
   assign mem[453759:453728] = 32'b00000111000110101110111011001000;
   assign mem[453791:453760] = 32'b00000010111000000010010010101000;
   assign mem[453823:453792] = 32'b00001000011110010110111100000000;
   assign mem[453855:453824] = 32'b11111100010011011000101110111000;
   assign mem[453887:453856] = 32'b00000000010011101000011001010010;
   assign mem[453919:453888] = 32'b11111100000000000101011000100100;
   assign mem[453951:453920] = 32'b00000001011000010100101011110000;
   assign mem[453983:453952] = 32'b00000010001000100111010110101000;
   assign mem[454015:453984] = 32'b11110111101110111010100011100000;
   assign mem[454047:454016] = 32'b00000001001101000011001011110010;
   assign mem[454079:454048] = 32'b00000011110000000001010100101000;
   assign mem[454111:454080] = 32'b00000110111100101011111001111000;
   assign mem[454143:454112] = 32'b11111010000010000011100110001000;
   assign mem[454175:454144] = 32'b11111111101011101101000011100011;
   assign mem[454207:454176] = 32'b11111011001111101001011011011000;
   assign mem[454239:454208] = 32'b11111010000000000101100000100000;
   assign mem[454271:454240] = 32'b00000001000110001010101101101010;
   assign mem[454303:454272] = 32'b00000011101010101001111100110100;
   assign mem[454335:454304] = 32'b11111010101111001010010100010000;
   assign mem[454367:454336] = 32'b00000010101101111010111011011000;
   assign mem[454399:454368] = 32'b00000000110110001000111011111111;
   assign mem[454431:454400] = 32'b00000001011110001110011110111100;
   assign mem[454463:454432] = 32'b00000100100010010001101000001000;
   assign mem[454495:454464] = 32'b00000100110000111111001011101000;
   assign mem[454527:454496] = 32'b11110111000101111110110000110000;
   assign mem[454559:454528] = 32'b00000110011010001001110100110000;
   assign mem[454591:454560] = 32'b11111110110111001111010100110100;
   assign mem[454623:454592] = 32'b11111001001101100111001001010000;
   assign mem[454655:454624] = 32'b11111001110100100100111110010000;
   assign mem[454687:454656] = 32'b11111111000010101101010010010101;
   assign mem[454719:454688] = 32'b00000011010100100011100010111100;
   assign mem[454751:454720] = 32'b00000101010010100001111110101000;
   assign mem[454783:454752] = 32'b11111001100001001011000010010000;
   assign mem[454815:454784] = 32'b00000000111001110001010100100010;
   assign mem[454847:454816] = 32'b00000000010010110001101010011111;
   assign mem[454879:454848] = 32'b11111011001101010000100000111000;
   assign mem[454911:454880] = 32'b00000110001110010010100100101000;
   assign mem[454943:454912] = 32'b00000010101001110100101001010100;
   assign mem[454975:454944] = 32'b11111000101101010110011101100000;
   assign mem[455007:454976] = 32'b00000001011010010100100100010110;
   assign mem[455039:455008] = 32'b11111110110110111001010001110100;
   assign mem[455071:455040] = 32'b00000011100110111000111001111000;
   assign mem[455103:455072] = 32'b11111101101000110111101101010100;
   assign mem[455135:455104] = 32'b00001000010111010010011000110000;
   assign mem[455167:455136] = 32'b11111101111001010100100010110100;
   assign mem[455199:455168] = 32'b11111011001111100000101001100000;
   assign mem[455231:455200] = 32'b11111111001010011010000111000001;
   assign mem[455263:455232] = 32'b00000010101010111111011101001100;
   assign mem[455295:455264] = 32'b11111100001000100011110001011000;
   assign mem[455327:455296] = 32'b00000111000000011001001110101000;
   assign mem[455359:455328] = 32'b11111000010110100000100110000000;
   assign mem[455391:455360] = 32'b11110110101010010100010000110000;
   assign mem[455423:455392] = 32'b00000101001011001000010110011000;
   assign mem[455455:455424] = 32'b11110111000110101011011000110000;
   assign mem[455487:455456] = 32'b00000100111110011110111101011000;
   assign mem[455519:455488] = 32'b00000011011110101010011000010000;
   assign mem[455551:455520] = 32'b00000010110011111101000010011000;
   assign mem[455583:455552] = 32'b11101111101100000101010101100000;
   assign mem[455615:455584] = 32'b00000101000001100101010111000000;
   assign mem[455647:455616] = 32'b11111001000111101110011001001000;
   assign mem[455679:455648] = 32'b00000100010100000111001111011000;
   assign mem[455711:455680] = 32'b00000101001001011001011011101000;
   assign mem[455743:455712] = 32'b00000000110011001101010010011101;
   assign mem[455775:455744] = 32'b00000101001111011110011101100000;
   assign mem[455807:455776] = 32'b00000000110010010010110001001100;
   assign mem[455839:455808] = 32'b11111011111001110011110111011000;
   assign mem[455871:455840] = 32'b00000001111010011001100000101100;
   assign mem[455903:455872] = 32'b00000011110111010011010110000100;
   assign mem[455935:455904] = 32'b11110100001100010001011001000000;
   assign mem[455967:455936] = 32'b00000010010111011101010101001100;
   assign mem[455999:455968] = 32'b11111100011001001000000000010100;
   assign mem[456031:456000] = 32'b11111100000110001010100101100100;
   assign mem[456063:456032] = 32'b00001001110000110110100011000000;
   assign mem[456095:456064] = 32'b00000010101101010000101000010100;
   assign mem[456127:456096] = 32'b11111000010100011000111001101000;
   assign mem[456159:456128] = 32'b00000000100011110101111101010111;
   assign mem[456191:456160] = 32'b11111111100000110011101000001100;
   assign mem[456223:456192] = 32'b00000101100001100111100010100000;
   assign mem[456255:456224] = 32'b11111100101011000100000110111000;
   assign mem[456287:456256] = 32'b00000001001011011110111111101110;
   assign mem[456319:456288] = 32'b11111111001000111111110101000100;
   assign mem[456351:456320] = 32'b00000010111100111111001000011100;
   assign mem[456383:456352] = 32'b00001100111001001011011000100000;
   assign mem[456415:456384] = 32'b00000101100110001111010000010000;
   assign mem[456447:456416] = 32'b11111100110011110100110101101000;
   assign mem[456479:456448] = 32'b11111010011011100011111010100000;
   assign mem[456511:456480] = 32'b11111110111100001000000110000000;
   assign mem[456543:456512] = 32'b11111101011010111100001000011100;
   assign mem[456575:456544] = 32'b11110000000011001000110011000000;
   assign mem[456607:456576] = 32'b11111100101100111101000101101000;
   assign mem[456639:456608] = 32'b11111011101101010000001111011000;
   assign mem[456671:456640] = 32'b11110110111000111010011110010000;
   assign mem[456703:456672] = 32'b11110010100000011001011111010000;
   assign mem[456735:456704] = 32'b00000111000001001011111110101000;
   assign mem[456767:456736] = 32'b00001001110001010110110010010000;
   assign mem[456799:456768] = 32'b11110111110110110010100000010000;
   assign mem[456831:456800] = 32'b00000000011010011001001100000111;
   assign mem[456863:456832] = 32'b11110101010111101010010001000000;
   assign mem[456895:456864] = 32'b11101110001000010000101000100000;
   assign mem[456927:456896] = 32'b00000010001000010010111100101000;
   assign mem[456959:456928] = 32'b00000000100001110001111101111110;
   assign mem[456991:456960] = 32'b11101100000011101111000000100000;
   assign mem[457023:456992] = 32'b00000110101101101011010111101000;
   assign mem[457055:457024] = 32'b11111100000011011100010011110000;
   assign mem[457087:457056] = 32'b11110100010110010010000100010000;
   assign mem[457119:457088] = 32'b00000110010001101110111010100000;
   assign mem[457151:457120] = 32'b11110001110000010011011111100000;
   assign mem[457183:457152] = 32'b11110010100111001001010000110000;
   assign mem[457215:457184] = 32'b00000100010000101100000111010000;
   assign mem[457247:457216] = 32'b00000010110100011110000000110100;
   assign mem[457279:457248] = 32'b00000110000101000101101101011000;
   assign mem[457311:457280] = 32'b00000000011110100010010000110011;
   assign mem[457343:457312] = 32'b11111110010111111111100101001110;
   assign mem[457375:457344] = 32'b00000001111110010110100110111010;
   assign mem[457407:457376] = 32'b00000101011000010000010001101000;
   assign mem[457439:457408] = 32'b11111000100100110110101111011000;
   assign mem[457471:457440] = 32'b00000100101101000011100101010000;
   assign mem[457503:457472] = 32'b11111110111110010000110101110000;
   assign mem[457535:457504] = 32'b11100011000111101111110111000000;
   assign mem[457567:457536] = 32'b00000001100100001011100111011010;
   assign mem[457599:457568] = 32'b11111100111011110111100000101100;
   assign mem[457631:457600] = 32'b00000111000011100000001110010000;
   assign mem[457663:457632] = 32'b11110110010011000101000100110000;
   assign mem[457695:457664] = 32'b11111001010110100000001101001000;
   assign mem[457727:457696] = 32'b00001000001010010011111111000000;
   assign mem[457759:457728] = 32'b00000100010011100110001111010000;
   assign mem[457791:457760] = 32'b00000011001110010011111000000100;
   assign mem[457823:457792] = 32'b11111100010100001000001001010000;
   assign mem[457855:457824] = 32'b00000011110111010010100110000100;
   assign mem[457887:457856] = 32'b11111100010110111011101111100000;
   assign mem[457919:457888] = 32'b00000101011010001011001101011000;
   assign mem[457951:457920] = 32'b00000110101010111110001100001000;
   assign mem[457983:457952] = 32'b00000001010001000000101110000000;
   assign mem[458015:457984] = 32'b00000000111001010111010111000110;
   assign mem[458047:458016] = 32'b11111111001100010101101010001101;
   assign mem[458079:458048] = 32'b11111000000111000100000111100000;
   assign mem[458111:458080] = 32'b11111100001101101010001110111100;
   assign mem[458143:458112] = 32'b00000101100111110100111011101000;
   assign mem[458175:458144] = 32'b11111101111000101010111010000100;
   assign mem[458207:458176] = 32'b00000001101111001111000010110000;
   assign mem[458239:458208] = 32'b11111100110110101101111111011000;
   assign mem[458271:458240] = 32'b00001001110101100100011000100000;
   assign mem[458303:458272] = 32'b00000000001011011111010100111111;
   assign mem[458335:458304] = 32'b11111011100010000000000111100000;
   assign mem[458367:458336] = 32'b11111010100111001010011101111000;
   assign mem[458399:458368] = 32'b11111110111000100110010100011100;
   assign mem[458431:458400] = 32'b11111111000111100110011001001010;
   assign mem[458463:458432] = 32'b00000100000000110011111000110000;
   assign mem[458495:458464] = 32'b11111101111011101110001101100000;
   assign mem[458527:458496] = 32'b00000011001011101111110100100000;
   assign mem[458559:458528] = 32'b11111011101110001011101101110000;
   assign mem[458591:458560] = 32'b11110001101010001111100101010000;
   assign mem[458623:458592] = 32'b00001000101110101100000110000000;
   assign mem[458655:458624] = 32'b11110110100110000100000100110000;
   assign mem[458687:458656] = 32'b11110000000001000011000101110000;
   assign mem[458719:458688] = 32'b00000101101110011010110011110000;
   assign mem[458751:458720] = 32'b00001000010011011100000111100000;
   assign mem[458783:458752] = 32'b11101111111000011001110101100000;
   assign mem[458815:458784] = 32'b00000111100000101101101100010000;
   assign mem[458847:458816] = 32'b11111011001001010111010011010000;
   assign mem[458879:458848] = 32'b00000101111001001000000100111000;
   assign mem[458911:458880] = 32'b00000101101101100101110111000000;
   assign mem[458943:458912] = 32'b00000011001010001101100010000100;
   assign mem[458975:458944] = 32'b11111101010111001110010100110100;
   assign mem[459007:458976] = 32'b11100111110011011100010110000000;
   assign mem[459039:459008] = 32'b00000000100110001010001101101100;
   assign mem[459071:459040] = 32'b11111000001010100000101010011000;
   assign mem[459103:459072] = 32'b00000001001101001111101010100010;
   assign mem[459135:459104] = 32'b00000010110111010110010001100000;
   assign mem[459167:459136] = 32'b00000101101010000111101010100000;
   assign mem[459199:459168] = 32'b11111111010010111010100111011000;
   assign mem[459231:459200] = 32'b11111001101100010100001111111000;
   assign mem[459263:459232] = 32'b00001111110111100000111100110000;
   assign mem[459295:459264] = 32'b00000111110001111010001011100000;
   assign mem[459327:459296] = 32'b00001001011111010111110110110000;
   assign mem[459359:459328] = 32'b11110100101001110011110111110000;
   assign mem[459391:459360] = 32'b00000111000111011001101101110000;
   assign mem[459423:459392] = 32'b11101101101101000001010001000000;
   assign mem[459455:459424] = 32'b00000011010001111011011111000100;
   assign mem[459487:459456] = 32'b11110110001001111100000110100000;
   assign mem[459519:459488] = 32'b11111101011000111110110101000000;
   assign mem[459551:459520] = 32'b00000100101101110011101011001000;
   assign mem[459583:459552] = 32'b11111000100111110110001011100000;
   assign mem[459615:459584] = 32'b00000010000010011011100001011000;
   assign mem[459647:459616] = 32'b00000001110100011111111011000010;
   assign mem[459679:459648] = 32'b11111011010110001111111110100000;
   assign mem[459711:459680] = 32'b00000000000111110010001111011010;
   assign mem[459743:459712] = 32'b00000010111100001101111011101100;
   assign mem[459775:459744] = 32'b11111001010011001000010100100000;
   assign mem[459807:459776] = 32'b00000101010010100001101111001000;
   assign mem[459839:459808] = 32'b11111100001010010101111101001100;
   assign mem[459871:459840] = 32'b11111101111000011011100000111000;
   assign mem[459903:459872] = 32'b00001000010111100111110101110000;
   assign mem[459935:459904] = 32'b11110110001010000010111111000000;
   assign mem[459967:459936] = 32'b00000000011110100111010001100001;
   assign mem[459999:459968] = 32'b11110001101101001010001100100000;
   assign mem[460031:460000] = 32'b00000011100001000111001100011000;
   assign mem[460063:460032] = 32'b11111100110010100011000111011100;
   assign mem[460095:460064] = 32'b11111100010101100101011101001100;
   assign mem[460127:460096] = 32'b11111010011111011011111010111000;
   assign mem[460159:460128] = 32'b11111111110010011010110011010011;
   assign mem[460191:460160] = 32'b11110100101101100101001111000000;
   assign mem[460223:460192] = 32'b00001010001010110011011100010000;
   assign mem[460255:460224] = 32'b11110110001110000010000000100000;
   assign mem[460287:460256] = 32'b11111101101001110110110101000100;
   assign mem[460319:460288] = 32'b00000101000011010000011101110000;
   assign mem[460351:460320] = 32'b11111100010110101011000001001000;
   assign mem[460383:460352] = 32'b11110110001000100110000101000000;
   assign mem[460415:460384] = 32'b00000100100101011001110011111000;
   assign mem[460447:460416] = 32'b00000000001111010111111010001101;
   assign mem[460479:460448] = 32'b00000111110111100100110001011000;
   assign mem[460511:460480] = 32'b00000001100010011000011111001010;
   assign mem[460543:460512] = 32'b11111111100111001010101101111101;
   assign mem[460575:460544] = 32'b11111100100000000001001111010000;
   assign mem[460607:460576] = 32'b00000000101010010011001110100100;
   assign mem[460639:460608] = 32'b11111110100010011011111110111000;
   assign mem[460671:460640] = 32'b11111101110100001101100111001000;
   assign mem[460703:460672] = 32'b00000000001011000111111111011001;
   assign mem[460735:460704] = 32'b11111011101110110010001101001000;
   assign mem[460767:460736] = 32'b11111111101000111010010100010110;
   assign mem[460799:460768] = 32'b00000001100001100110001110011110;
   assign mem[460831:460800] = 32'b00000100110111101111111010100000;
   assign mem[460863:460832] = 32'b00000001110110000011011010011100;
   assign mem[460895:460864] = 32'b00000010001110111011100011111000;
   assign mem[460927:460896] = 32'b00000111001000110101101011011000;
   assign mem[460959:460928] = 32'b11111101100101001001111010010100;
   assign mem[460991:460960] = 32'b00000011010111000010101010111000;
   assign mem[461023:460992] = 32'b11111010101101111001001001100000;
   assign mem[461055:461024] = 32'b11111011000001110011101110110000;
   assign mem[461087:461056] = 32'b11110010111110000011100101110000;
   assign mem[461119:461088] = 32'b11111111110000101111011111110101;
   assign mem[461151:461120] = 32'b11111100100011010100000110111000;
   assign mem[461183:461152] = 32'b00000010010000001010010111111000;
   assign mem[461215:461184] = 32'b11111000110110001011011111111000;
   assign mem[461247:461216] = 32'b00000001001011011001110100100110;
   assign mem[461279:461248] = 32'b00000100000000000110000111011000;
   assign mem[461311:461280] = 32'b11111010100010010111000010101000;
   assign mem[461343:461312] = 32'b11110110101101001011010000110000;
   assign mem[461375:461344] = 32'b00000101101000000010111011010000;
   assign mem[461407:461376] = 32'b11110110111000010101100011100000;
   assign mem[461439:461408] = 32'b00000100100000110110100110001000;
   assign mem[461471:461440] = 32'b00000001010100101001100010001100;
   assign mem[461503:461472] = 32'b00000011010110101001001010110000;
   assign mem[461535:461504] = 32'b00000000111100000010101101000100;
   assign mem[461567:461536] = 32'b11111101111011000101101101100000;
   assign mem[461599:461568] = 32'b11111000010000101111101011000000;
   assign mem[461631:461600] = 32'b00000000001101111001000100010110;
   assign mem[461663:461632] = 32'b00000011010001000001111100000000;
   assign mem[461695:461664] = 32'b11111101011110010010110010010000;
   assign mem[461727:461696] = 32'b11111111100001000101010010101101;
   assign mem[461759:461728] = 32'b11111100001011001010110001010000;
   assign mem[461791:461760] = 32'b11111100001011101010110111100000;
   assign mem[461823:461792] = 32'b00001000100001011000001100000000;
   assign mem[461855:461824] = 32'b11111010000000101101100110011000;
   assign mem[461887:461856] = 32'b11110111000110000010110111100000;
   assign mem[461919:461888] = 32'b11111110000110110101001110001010;
   assign mem[461951:461920] = 32'b00001100100111010101011010110000;
   assign mem[461983:461952] = 32'b11110110101011000001011101010000;
   assign mem[462015:461984] = 32'b00000011101101101100110110100100;
   assign mem[462047:462016] = 32'b11111111100101001110010001011110;
   assign mem[462079:462048] = 32'b00000011000111100010000001101100;
   assign mem[462111:462080] = 32'b00001000100000010001110110010000;
   assign mem[462143:462112] = 32'b11110111010101101101101000010000;
   assign mem[462175:462144] = 32'b00000011010001010101111000010100;
   assign mem[462207:462176] = 32'b00000100011100111000001000100000;
   assign mem[462239:462208] = 32'b11111000110011001110001010011000;
   assign mem[462271:462240] = 32'b00000011011011001101010110000100;
   assign mem[462303:462272] = 32'b00000100110101011011001001000000;
   assign mem[462335:462304] = 32'b11101011011110111000101100000000;
   assign mem[462367:462336] = 32'b11111101100010101100000001010000;
   assign mem[462399:462368] = 32'b11111111001000110001111111010001;
   assign mem[462431:462400] = 32'b00000001011111110001110010000100;
   assign mem[462463:462432] = 32'b00001000010010011001111101100000;
   assign mem[462495:462464] = 32'b11111111001000101100101110110011;
   assign mem[462527:462496] = 32'b11111111110100101010101001100100;
   assign mem[462559:462528] = 32'b11110101100001001101110111000000;
   assign mem[462591:462560] = 32'b00000001100110111010111111010010;
   assign mem[462623:462592] = 32'b00000000010011111101011001110101;
   assign mem[462655:462624] = 32'b11110111110110110101011000010000;
   assign mem[462687:462656] = 32'b00000111010001110101010010001000;
   assign mem[462719:462688] = 32'b00000001001011100011111110110000;
   assign mem[462751:462720] = 32'b00001000001011010001001010100000;
   assign mem[462783:462752] = 32'b00000000100101010011010110110110;
   assign mem[462815:462784] = 32'b00000111010001000101011110110000;
   assign mem[462847:462816] = 32'b11111111100010110100001011110010;
   assign mem[462879:462848] = 32'b11111000111110111000001000111000;
   assign mem[462911:462880] = 32'b11111111001101010100111110000001;
   assign mem[462943:462912] = 32'b00000101001010101100100011000000;
   assign mem[462975:462944] = 32'b11111000010110001101100110011000;
   assign mem[463007:462976] = 32'b00000010000110010101110100101000;
   assign mem[463039:463008] = 32'b11110011001101011000010001010000;
   assign mem[463071:463040] = 32'b00000010001011000010110011101100;
   assign mem[463103:463072] = 32'b11110100110110011111011110110000;
   assign mem[463135:463104] = 32'b00000011001101100100001110101100;
   assign mem[463167:463136] = 32'b00001100111000101101111001000000;
   assign mem[463199:463168] = 32'b11110111111110110111000011100000;
   assign mem[463231:463200] = 32'b00001000101010001011100010100000;
   assign mem[463263:463232] = 32'b11111011001010101001000011110000;
   assign mem[463295:463264] = 32'b11110111100001100101001001110000;
   assign mem[463327:463296] = 32'b11101111011010111010010100000000;
   assign mem[463359:463328] = 32'b11111111101001111011101111100111;
   assign mem[463391:463360] = 32'b00000101101011010000111001101000;
   assign mem[463423:463392] = 32'b00000001101010010111010100111100;
   assign mem[463455:463424] = 32'b00000111000011100010101010110000;
   assign mem[463487:463456] = 32'b11111111001010011101101110000001;
   assign mem[463519:463488] = 32'b11110110000111100100110111010000;
   assign mem[463551:463520] = 32'b11111100101010101000000011011100;
   assign mem[463583:463552] = 32'b00000111101010001111111100011000;
   assign mem[463615:463584] = 32'b11110111100110001001111000000000;
   assign mem[463647:463616] = 32'b11111110101011110000100001001100;
   assign mem[463679:463648] = 32'b11111011110100001010111111101000;
   assign mem[463711:463680] = 32'b00000010100110000011101000111000;
   assign mem[463743:463712] = 32'b11111111101010000100001000111101;
   assign mem[463775:463744] = 32'b00000000101011100000000000100111;
   assign mem[463807:463776] = 32'b11111101101010001100101111011100;
   assign mem[463839:463808] = 32'b11111111010001001110011110010011;
   assign mem[463871:463840] = 32'b00000010110001110110100111110100;
   assign mem[463903:463872] = 32'b00000100001110110101010010101000;
   assign mem[463935:463904] = 32'b11110111111001100100010100110000;
   assign mem[463967:463936] = 32'b11111101111110010100111100110100;
   assign mem[463999:463968] = 32'b11111111100100111101111000110010;
   assign mem[464031:464000] = 32'b00000010011010000101111101101000;
   assign mem[464063:464032] = 32'b00000001010111000011110111000110;
   assign mem[464095:464064] = 32'b00000100100100101011011001010000;
   assign mem[464127:464096] = 32'b00000001100101011100110000111100;
   assign mem[464159:464128] = 32'b11111011010001001110111111011000;
   assign mem[464191:464160] = 32'b11111101110110101000111100101100;
   assign mem[464223:464192] = 32'b00000010111001001110011010011000;
   assign mem[464255:464224] = 32'b11111000001000001001011010110000;
   assign mem[464287:464256] = 32'b00000000010100001001101011110001;
   assign mem[464319:464288] = 32'b11111001010011111001000111111000;
   assign mem[464351:464320] = 32'b00010001110100001010001001000000;
   assign mem[464383:464352] = 32'b00000101111100110101000100010000;
   assign mem[464415:464384] = 32'b00000000001000010110000011001110;
   assign mem[464447:464416] = 32'b11111100110000110010001111111100;
   assign mem[464479:464448] = 32'b11110111010101111101110110010000;
   assign mem[464511:464480] = 32'b11111111100110101001010110000001;
   assign mem[464543:464512] = 32'b00000100111010111010011001101000;
   assign mem[464575:464544] = 32'b00000000111101111110101101110001;
   assign mem[464607:464576] = 32'b00000001100101001111110000101110;
   assign mem[464639:464608] = 32'b11110001110011000110101001100000;
   assign mem[464671:464640] = 32'b00001001010001111100111110110000;
   assign mem[464703:464672] = 32'b00000100100000111110111011111000;
   assign mem[464735:464704] = 32'b00000110001100100010011010100000;
   assign mem[464767:464736] = 32'b11111110000111001011100001000100;
   assign mem[464799:464768] = 32'b11110100011011010100011001010000;
   assign mem[464831:464800] = 32'b11111101011000010110011110000000;
   assign mem[464863:464832] = 32'b00000110010010100001011100111000;
   assign mem[464895:464864] = 32'b11111101101110011100011100100100;
   assign mem[464927:464896] = 32'b00000110000010101111000110110000;
   assign mem[464959:464928] = 32'b11101101111010000100111001000000;
   assign mem[464991:464960] = 32'b00000001110100011000111110011010;
   assign mem[465023:464992] = 32'b11111010100001101100010100010000;
   assign mem[465055:465024] = 32'b11111010101100111100111000010000;
   assign mem[465087:465056] = 32'b00000111001001010010101000110000;
   assign mem[465119:465088] = 32'b00000011100111001000011100001100;
   assign mem[465151:465120] = 32'b00001000011101110111101000010000;
   assign mem[465183:465152] = 32'b00000101000010010100011010110000;
   assign mem[465215:465184] = 32'b00000001101101001010101010010010;
   assign mem[465247:465216] = 32'b11110101111100101011010110110000;
   assign mem[465279:465248] = 32'b11111000100100110101100110100000;
   assign mem[465311:465280] = 32'b11110100111100011100010100110000;
   assign mem[465343:465312] = 32'b00001011011101101000101100000000;
   assign mem[465375:465344] = 32'b11110011110101111001110101100000;
   assign mem[465407:465376] = 32'b11110101110100101000000001010000;
   assign mem[465439:465408] = 32'b00000111111011000011100001111000;
   assign mem[465471:465440] = 32'b11110111111100111100000011110000;
   assign mem[465503:465472] = 32'b11110111101010101010000110000000;
   assign mem[465535:465504] = 32'b00001100101100111101101100110000;
   assign mem[465567:465536] = 32'b11110100010101111111100110010000;
   assign mem[465599:465568] = 32'b00001010110111011011010110010000;
   assign mem[465631:465600] = 32'b00000001000001101110101000001100;
   assign mem[465663:465632] = 32'b11111101101100010011001111110000;
   assign mem[465695:465664] = 32'b11111111110101100100111011100010;
   assign mem[465727:465696] = 32'b11111101101110101000111100010000;
   assign mem[465759:465728] = 32'b00000011101000100000010010110100;
   assign mem[465791:465760] = 32'b11111101111000101000100101110000;
   assign mem[465823:465792] = 32'b11111100001100101010010000111000;
   assign mem[465855:465824] = 32'b00000011100010010100011111000000;
   assign mem[465887:465856] = 32'b00000010111001001000110100001000;
   assign mem[465919:465888] = 32'b11111100100000111110100011111100;
   assign mem[465951:465920] = 32'b00000000110110100110001110100000;
   assign mem[465983:465952] = 32'b00000000011011000001101010100100;
   assign mem[466015:465984] = 32'b00000110000001101101011000100000;
   assign mem[466047:466016] = 32'b00000001000010111010011000100100;
   assign mem[466079:466048] = 32'b11111101000000001101010001000100;
   assign mem[466111:466080] = 32'b00000110000001010110001110101000;
   assign mem[466143:466112] = 32'b00000010001010000001101011000000;
   assign mem[466175:466144] = 32'b11111011101100011110100011101000;
   assign mem[466207:466176] = 32'b11111110111110100000001001111000;
   assign mem[466239:466208] = 32'b11110101100010110111001001000000;
   assign mem[466271:466240] = 32'b11111111011101110000111001000111;
   assign mem[466303:466272] = 32'b00000001000011101110011100010110;
   assign mem[466335:466304] = 32'b00000010001000111100101101010100;
   assign mem[466367:466336] = 32'b00000010111000101111011011101000;
   assign mem[466399:466368] = 32'b11111100011000000000100100001100;
   assign mem[466431:466400] = 32'b00000010111000000011010001110100;
   assign mem[466463:466432] = 32'b11111011100011011110111100100000;
   assign mem[466495:466464] = 32'b11111111010011000000111001100111;
   assign mem[466527:466496] = 32'b11111000001110100000111110111000;
   assign mem[466559:466528] = 32'b00000000000010110000101001001101;
   assign mem[466591:466560] = 32'b00000010010111111011010100000100;
   assign mem[466623:466592] = 32'b11101011100111001100110011000000;
   assign mem[466655:466624] = 32'b00000001011111101110001010100100;
   assign mem[466687:466656] = 32'b00001000001010111000101000100000;
   assign mem[466719:466688] = 32'b11111101101001100110001000011100;
   assign mem[466751:466720] = 32'b00000110001111011011100110100000;
   assign mem[466783:466752] = 32'b11111111000001111110110100100110;
   assign mem[466815:466784] = 32'b11111101001100011011110010110000;
   assign mem[466847:466816] = 32'b00000111001100100111010000101000;
   assign mem[466879:466848] = 32'b11111101001101010100001110010000;
   assign mem[466911:466880] = 32'b11011111011001101010100111000000;
   assign mem[466943:466912] = 32'b00000111111001110001010011001000;
   assign mem[466975:466944] = 32'b11111001001110001100011010011000;
   assign mem[467007:466976] = 32'b11110110011110000001000010110000;
   assign mem[467039:467008] = 32'b00000111010110100000101110000000;
   assign mem[467071:467040] = 32'b11110101011001011111110100010000;
   assign mem[467103:467072] = 32'b11110110001000010111111000010000;
   assign mem[467135:467104] = 32'b00000110011010110101110011011000;
   assign mem[467167:467136] = 32'b11111100000111101011110011001100;
   assign mem[467199:467168] = 32'b00001000100001110100110110100000;
   assign mem[467231:467200] = 32'b11111111111011110000110001100001;
   assign mem[467263:467232] = 32'b00000000101110010000010000001011;
   assign mem[467295:467264] = 32'b11111100101101000111001011011000;
   assign mem[467327:467296] = 32'b11111101100111100111010010011100;
   assign mem[467359:467328] = 32'b11111000110111010011001100100000;
   assign mem[467391:467360] = 32'b11111111110110111111110110010011;
   assign mem[467423:467392] = 32'b00000001101110110110100010001110;
   assign mem[467455:467424] = 32'b11111001001110111010010011011000;
   assign mem[467487:467456] = 32'b00000001101010010011111011111100;
   assign mem[467519:467488] = 32'b11111011101100001101010110111000;
   assign mem[467551:467520] = 32'b11111110100111100011000111111000;
   assign mem[467583:467552] = 32'b00000101000101010111110100010000;
   assign mem[467615:467584] = 32'b00000001100000010000101111111100;
   assign mem[467647:467616] = 32'b00000001000101011110110101101100;
   assign mem[467679:467648] = 32'b11111000111100101010011100100000;
   assign mem[467711:467680] = 32'b11111111110100111100000100100001;
   assign mem[467743:467712] = 32'b00000010101110100000100100000100;
   assign mem[467775:467744] = 32'b11110011010100111110010111000000;
   assign mem[467807:467776] = 32'b00000000000010110111100010000101;
   assign mem[467839:467808] = 32'b11111101100100000100011111000100;
   assign mem[467871:467840] = 32'b00000011010011101110000010011000;
   assign mem[467903:467872] = 32'b00000010010011011011101011010100;
   assign mem[467935:467904] = 32'b11111101100110010101110100001100;
   assign mem[467967:467936] = 32'b00000000101001011100101001101111;
   assign mem[467999:467968] = 32'b11111011110100000101011101111000;
   assign mem[468031:468000] = 32'b00000001011111110110000010011100;
   assign mem[468063:468032] = 32'b00000010000001001000111001010000;
   assign mem[468095:468064] = 32'b11111011000110000001101010000000;
   assign mem[468127:468096] = 32'b11111100100100001100000101011000;
   assign mem[468159:468128] = 32'b11111010101110100010100000110000;
   assign mem[468191:468160] = 32'b11111010110010100110011011111000;
   assign mem[468223:468192] = 32'b00000010100011010000001011111100;
   assign mem[468255:468224] = 32'b11110011110000101100111001100000;
   assign mem[468287:468256] = 32'b11101100111010011111000000000000;
   assign mem[468319:468288] = 32'b00000100010100000010001100111000;
   assign mem[468351:468320] = 32'b00000000010111010000011001010011;
   assign mem[468383:468352] = 32'b11110000010101000011111010000000;
   assign mem[468415:468384] = 32'b00000110100101001000010110001000;
   assign mem[468447:468416] = 32'b00000000100011011001010000110101;
   assign mem[468479:468448] = 32'b00000110000110110110010011000000;
   assign mem[468511:468480] = 32'b11111001101111000010001011010000;
   assign mem[468543:468512] = 32'b00000100011110101000111011010000;
   assign mem[468575:468544] = 32'b11110110111100101001011000010000;
   assign mem[468607:468576] = 32'b00000001111110011110111111001000;
   assign mem[468639:468608] = 32'b11111001000010001000011100011000;
   assign mem[468671:468640] = 32'b00001111000001011011000001110000;
   assign mem[468703:468672] = 32'b00000000101001010000000010100000;
   assign mem[468735:468704] = 32'b11111011011101101111100001000000;
   assign mem[468767:468736] = 32'b00000101000010011111000100011000;
   assign mem[468799:468768] = 32'b11110110111010001011111110000000;
   assign mem[468831:468800] = 32'b00000010110010111101000001011000;
   assign mem[468863:468832] = 32'b11111001111110111111000101011000;
   assign mem[468895:468864] = 32'b11111111000110011111101111101011;
   assign mem[468927:468896] = 32'b11111101100111101001111111111000;
   assign mem[468959:468928] = 32'b00000010101001100100100110110100;
   assign mem[468991:468960] = 32'b00000011001000001100111111010000;
   assign mem[469023:468992] = 32'b00000011010111010111100111000000;
   assign mem[469055:469024] = 32'b11111010111010100110101001100000;
   assign mem[469087:469056] = 32'b11111110011111011001010110000110;
   assign mem[469119:469088] = 32'b11111111101010001100011010100001;
   assign mem[469151:469120] = 32'b00001011100100101110000011000000;
   assign mem[469183:469152] = 32'b11110110100010001101111011110000;
   assign mem[469215:469184] = 32'b11110111100100111000000011010000;
   assign mem[469247:469216] = 32'b00000110111110011100001001100000;
   assign mem[469279:469248] = 32'b11101100110010011011000000100000;
   assign mem[469311:469280] = 32'b00001010010010001010010111010000;
   assign mem[469343:469312] = 32'b11111011101101000000100001100000;
   assign mem[469375:469344] = 32'b11110001001011111010011010000000;
   assign mem[469407:469376] = 32'b11110101101100000010101111110000;
   assign mem[469439:469408] = 32'b00000100110011100101011100001000;
   assign mem[469471:469440] = 32'b00000100110011100111110100000000;
   assign mem[469503:469472] = 32'b00000010010110111001101110100000;
   assign mem[469535:469504] = 32'b11111001101001101011010101111000;
   assign mem[469567:469536] = 32'b00001010001001101010101111000000;
   assign mem[469599:469568] = 32'b11101100001001110111010100000000;
   assign mem[469631:469600] = 32'b00000111100101111011010101100000;
   assign mem[469663:469632] = 32'b00000001100000011111100101010110;
   assign mem[469695:469664] = 32'b11110101111000101111111111100000;
   assign mem[469727:469696] = 32'b11111111100111010100000010010111;
   assign mem[469759:469728] = 32'b11110101111001110100000001000000;
   assign mem[469791:469760] = 32'b11110100100100100111100010010000;
   assign mem[469823:469792] = 32'b00001010110011001001001110110000;
   assign mem[469855:469824] = 32'b00000001011000111000110001000100;
   assign mem[469887:469856] = 32'b00010001000011011001101110000000;
   assign mem[469919:469888] = 32'b11110100110111000110001001110000;
   assign mem[469951:469920] = 32'b00000111101010000110101010001000;
   assign mem[469983:469952] = 32'b11100111111101101000101100000000;
   assign mem[470015:469984] = 32'b11111010000000110111010101100000;
   assign mem[470047:470016] = 32'b11101110100010111100000100000000;
   assign mem[470079:470048] = 32'b00000100101101011111111011100000;
   assign mem[470111:470080] = 32'b11111100111000000010111001101100;
   assign mem[470143:470112] = 32'b00000010001010011001001101100100;
   assign mem[470175:470144] = 32'b00000110010011101010000110101000;
   assign mem[470207:470176] = 32'b00000010011001011100011110111100;
   assign mem[470239:470208] = 32'b11111111100100101000000010101000;
   assign mem[470271:470240] = 32'b11111110110101110100101111001010;
   assign mem[470303:470272] = 32'b11111101011000001110010110010000;
   assign mem[470335:470304] = 32'b00000000101010101101000010111110;
   assign mem[470367:470336] = 32'b11110110011011010001111000110000;
   assign mem[470399:470368] = 32'b00000001110000100110010001100000;
   assign mem[470431:470400] = 32'b11111100010110000100111100110100;
   assign mem[470463:470432] = 32'b00000100000001001010011100101000;
   assign mem[470495:470464] = 32'b00000001000111011001100101000000;
   assign mem[470527:470496] = 32'b11110010110111011101001111000000;
   assign mem[470559:470528] = 32'b00000000001010011010011100101001;
   assign mem[470591:470560] = 32'b11101110010011100000010101000000;
   assign mem[470623:470592] = 32'b11110000110010001001011000100000;
   assign mem[470655:470624] = 32'b00000000011010010000000011001110;
   assign mem[470687:470656] = 32'b11111111000111100101101110110000;
   assign mem[470719:470688] = 32'b00000001010110111100010110111000;
   assign mem[470751:470720] = 32'b11111010101001100111001110001000;
   assign mem[470783:470752] = 32'b11111110001001111010001011110000;
   assign mem[470815:470784] = 32'b11111101110000111110010110001000;
   assign mem[470847:470816] = 32'b11111100100111010011011011111000;
   assign mem[470879:470848] = 32'b00000010001011000001110001111100;
   assign mem[470911:470880] = 32'b11111100011010001111111111110000;
   assign mem[470943:470912] = 32'b11101011101101000010001000000000;
   assign mem[470975:470944] = 32'b00000010110000110101101111011000;
   assign mem[471007:470976] = 32'b11111011100010101101001011010000;
   assign mem[471039:471008] = 32'b00000101100010111010000100100000;
   assign mem[471071:471040] = 32'b00000001100010110011010011111010;
   assign mem[471103:471072] = 32'b11101000010100011001000111100000;
   assign mem[471135:471104] = 32'b00001011001010101000100111010000;
   assign mem[471167:471136] = 32'b00000100000101111010001110000000;
   assign mem[471199:471168] = 32'b11111100111011011010011110101100;
   assign mem[471231:471200] = 32'b11111100110010001000011010111100;
   assign mem[471263:471232] = 32'b00001000010100110000101111000000;
   assign mem[471295:471264] = 32'b11111000110110001101111011111000;
   assign mem[471327:471296] = 32'b00000011000100011011000110010100;
   assign mem[471359:471328] = 32'b11111101011000010000011101111100;
   assign mem[471391:471360] = 32'b11011111010100101110110101000000;
   assign mem[471423:471392] = 32'b00000111010000101000011101111000;
   assign mem[471455:471424] = 32'b11110010010100101001110100000000;
   assign mem[471487:471456] = 32'b00000111011001110111110011001000;
   assign mem[471519:471488] = 32'b11111000000111001101001011011000;
   assign mem[471551:471520] = 32'b00000111010110111111110100011000;
   assign mem[471583:471552] = 32'b11111011101100000011110011001000;
   assign mem[471615:471584] = 32'b00001000011000001111100111110000;
   assign mem[471647:471616] = 32'b00000010001011111100001111100000;
   assign mem[471679:471648] = 32'b11110111010100001100101100100000;
   assign mem[471711:471680] = 32'b11111100010000001110000010001100;
   assign mem[471743:471712] = 32'b00000010101100110101100100110100;
   assign mem[471775:471744] = 32'b00000111110000011110001011000000;
   assign mem[471807:471776] = 32'b00000101001110000011011010001000;
   assign mem[471839:471808] = 32'b11111010011010100001010100011000;
   assign mem[471871:471840] = 32'b11111010010010110101011100111000;
   assign mem[471903:471872] = 32'b00000001111101010101001001110010;
   assign mem[471935:471904] = 32'b11110100010111000111100111110000;
   assign mem[471967:471936] = 32'b00000001111100011110100101000110;
   assign mem[471999:471968] = 32'b11110110000110111010111001100000;
   assign mem[472031:472000] = 32'b00000001101010101110000000110000;
   assign mem[472063:472032] = 32'b00000011001111100011101001111100;
   assign mem[472095:472064] = 32'b11111110100101000001001101100010;
   assign mem[472127:472096] = 32'b11111101001011010100101111001100;
   assign mem[472159:472128] = 32'b11111110111101101011100110111100;
   assign mem[472191:472160] = 32'b11111100101100100100111111110100;
   assign mem[472223:472192] = 32'b00000001000101010110011110001010;
   assign mem[472255:472224] = 32'b11110101010010111110111000000000;
   assign mem[472287:472256] = 32'b11111110001101001110101111001110;
   assign mem[472319:472288] = 32'b11110110100010101010110011010000;
   assign mem[472351:472320] = 32'b00000010011010111110110101101000;
   assign mem[472383:472352] = 32'b00000010001000100111001011111000;
   assign mem[472415:472384] = 32'b00000100001011011000011100010000;
   assign mem[472447:472416] = 32'b11111011101100101000011110111000;
   assign mem[472479:472448] = 32'b11111011001001100010001000100000;
   assign mem[472511:472480] = 32'b11111011111011011110100111000000;
   assign mem[472543:472512] = 32'b00000100110101110010100001100000;
   assign mem[472575:472544] = 32'b11111110100110011010111111001000;
   assign mem[472607:472576] = 32'b00000000110100010011100101000000;
   assign mem[472639:472608] = 32'b11111100001101000010110110110100;
   assign mem[472671:472640] = 32'b00000100010101100001110010010000;
   assign mem[472703:472672] = 32'b11110011000001011110100000100000;
   assign mem[472735:472704] = 32'b11111111100111000011110111000100;
   assign mem[472767:472736] = 32'b00000001111001101111011111110000;
   assign mem[472799:472768] = 32'b11111101011001001010010101100000;
   assign mem[472831:472800] = 32'b00000011111101111011110000000000;
   assign mem[472863:472832] = 32'b11111110011000000100101011011000;
   assign mem[472895:472864] = 32'b11111101011000110000101100100100;
   assign mem[472927:472896] = 32'b00000010000001101011000011101000;
   assign mem[472959:472928] = 32'b11111111010011010100010010101010;
   assign mem[472991:472960] = 32'b00000000010101110111100011111100;
   assign mem[473023:472992] = 32'b00000001011101111000001010111100;
   assign mem[473055:473024] = 32'b11111000011001101111001101111000;
   assign mem[473087:473056] = 32'b11111111011010111001101011110110;
   assign mem[473119:473088] = 32'b11111111001010010111111010011000;
   assign mem[473151:473120] = 32'b00000001011111111110000010010110;
   assign mem[473183:473152] = 32'b00000001111011001000101000101110;
   assign mem[473215:473184] = 32'b11111110111100011110110001000000;
   assign mem[473247:473216] = 32'b00000000100011000101000101001000;
   assign mem[473279:473248] = 32'b11111111000111110011001011010010;
   assign mem[473311:473280] = 32'b00000100110010100101101110101000;
   assign mem[473343:473312] = 32'b11110001001011011010111100000000;
   assign mem[473375:473344] = 32'b00000001010000011000110001011100;
   assign mem[473407:473376] = 32'b00000001111100011001111001011000;
   assign mem[473439:473408] = 32'b11110110111010001100110111110000;
   assign mem[473471:473440] = 32'b00000100100111100011001101000000;
   assign mem[473503:473472] = 32'b00000010011011110000001111000100;
   assign mem[473535:473504] = 32'b11111010101011010111011101111000;
   assign mem[473567:473536] = 32'b00000011100001100110111011110100;
   assign mem[473599:473568] = 32'b00000000001110000010000100001100;
   assign mem[473631:473600] = 32'b00000101101101111001010001110000;
   assign mem[473663:473632] = 32'b00000000010110010001001010001100;
   assign mem[473695:473664] = 32'b00000100000111011000001001101000;
   assign mem[473727:473696] = 32'b00000001101101011111001010010000;
   assign mem[473759:473728] = 32'b11111010110111011001111001010000;
   assign mem[473791:473760] = 32'b00000001011111011110000010000000;
   assign mem[473823:473792] = 32'b00000010001101010000010101001000;
   assign mem[473855:473824] = 32'b11101101101001000101000001100000;
   assign mem[473887:473856] = 32'b11111100000101010111100111100000;
   assign mem[473919:473888] = 32'b11111110111011101000011010010000;
   assign mem[473951:473920] = 32'b11110111100011110110101111000000;
   assign mem[473983:473952] = 32'b00000010010010001100101010101100;
   assign mem[474015:473984] = 32'b11110000111010010000111001110000;
   assign mem[474047:474016] = 32'b00000011110110111000010011010100;
   assign mem[474079:474048] = 32'b11111110101110010010100101001100;
   assign mem[474111:474080] = 32'b00000000100010010111010101010100;
   assign mem[474143:474112] = 32'b11111010011010000110100100010000;
   assign mem[474175:474144] = 32'b00000010011100001000111000011100;
   assign mem[474207:474176] = 32'b11111101111000011110111110100000;
   assign mem[474239:474208] = 32'b00000110001101111000100101101000;
   assign mem[474271:474240] = 32'b00000000011101011101001001111011;
   assign mem[474303:474272] = 32'b00000100111111111000111001100000;
   assign mem[474335:474304] = 32'b11111101110011011010101001100100;
   assign mem[474367:474336] = 32'b00000001010011100010011010101010;
   assign mem[474399:474368] = 32'b11111110001101000110111110101010;
   assign mem[474431:474400] = 32'b00000000110011100000111001110010;
   assign mem[474463:474432] = 32'b11111110011000000011110111100000;
   assign mem[474495:474464] = 32'b11110110010100111111111111010000;
   assign mem[474527:474496] = 32'b11111111111010101010001001100101;
   assign mem[474559:474528] = 32'b00000001100101101100110010100010;
   assign mem[474591:474560] = 32'b00000000111111001001101000000100;
   assign mem[474623:474592] = 32'b00000000010010011110111010101000;
   assign mem[474655:474624] = 32'b00000101011100000100010001111000;
   assign mem[474687:474656] = 32'b00000010001000011010110100000000;
   assign mem[474719:474688] = 32'b00000010010000110011011010111000;
   assign mem[474751:474720] = 32'b11111000111110001101001100001000;
   assign mem[474783:474752] = 32'b00000001010101010010001110111010;
   assign mem[474815:474784] = 32'b11111011010100110101010000111000;
   assign mem[474847:474816] = 32'b11111110000010010111101000000000;
   assign mem[474879:474848] = 32'b11111101011010000100101100101000;
   assign mem[474911:474880] = 32'b11111111011000100110000110110000;
   assign mem[474943:474912] = 32'b11111111010000110111001000101010;
   assign mem[474975:474944] = 32'b00001110011011001110000001110000;
   assign mem[475007:474976] = 32'b11111010010001110101001011010000;
   assign mem[475039:475008] = 32'b11111110110011000101001011001010;
   assign mem[475071:475040] = 32'b11111110011111001000110010000110;
   assign mem[475103:475072] = 32'b00000011001100100100001111110100;
   assign mem[475135:475104] = 32'b00000000100100110010110110101011;
   assign mem[475167:475136] = 32'b11111011000101010111011011100000;
   assign mem[475199:475168] = 32'b00000101000001110100001101001000;
   assign mem[475231:475200] = 32'b11111101000111101111111111110100;
   assign mem[475263:475232] = 32'b00000111110100110111010001010000;
   assign mem[475295:475264] = 32'b00010011000011011110100010000000;
   assign mem[475327:475296] = 32'b00000000011000001100011111010110;
   assign mem[475359:475328] = 32'b11111110010100110000000110001100;
   assign mem[475391:475360] = 32'b11111110010110001101100111111100;
   assign mem[475423:475392] = 32'b11110110111100011011101010000000;
   assign mem[475455:475424] = 32'b11111001110000100001000001111000;
   assign mem[475487:475456] = 32'b11111101000000111010100000000100;
   assign mem[475519:475488] = 32'b11111001101001100010010111010000;
   assign mem[475551:475520] = 32'b00000000101001010101110111000001;
   assign mem[475583:475552] = 32'b00000010101000000011000101110100;
   assign mem[475615:475584] = 32'b00001010001000001001100011000000;
   assign mem[475647:475616] = 32'b11110111011001110000101011100000;
   assign mem[475679:475648] = 32'b11111010001001100010010101101000;
   assign mem[475711:475680] = 32'b11111100100010111011011001101100;
   assign mem[475743:475712] = 32'b00000100010110001010010011111000;
   assign mem[475775:475744] = 32'b11111000010001000111010001001000;
   assign mem[475807:475776] = 32'b00000100000101111101110101111000;
   assign mem[475839:475808] = 32'b11111000100010101010001110011000;
   assign mem[475871:475840] = 32'b11111001000010100010111011011000;
   assign mem[475903:475872] = 32'b11110101011100011011100000100000;
   assign mem[475935:475904] = 32'b11110001011010111100101100010000;
   assign mem[475967:475936] = 32'b00000111011110110100110001011000;
   assign mem[475999:475968] = 32'b00000000100100010110111010101101;
   assign mem[476031:476000] = 32'b11111111110000010100010110001111;
   assign mem[476063:476032] = 32'b11111000010001011010101100001000;
   assign mem[476095:476064] = 32'b00000001111110111011001110000010;
   assign mem[476127:476096] = 32'b00000000000111101011010100110010;
   assign mem[476159:476128] = 32'b00000000101111111111100110101110;
   assign mem[476191:476160] = 32'b00000010111001010100110000011000;
   assign mem[476223:476192] = 32'b00000001101110100100110010110000;
   assign mem[476255:476224] = 32'b00000000110010110001101110010000;
   assign mem[476287:476256] = 32'b11111111001010110010011100011011;
   assign mem[476319:476288] = 32'b11111001110101100000101110100000;
   assign mem[476351:476320] = 32'b11111011000101111100100111000000;
   assign mem[476383:476352] = 32'b00000001100111011100111110000100;
   assign mem[476415:476384] = 32'b11111010010101111011001111111000;
   assign mem[476447:476416] = 32'b11111101000110011011010011011100;
   assign mem[476479:476448] = 32'b11111100110001100010001010110000;
   assign mem[476511:476480] = 32'b11111000101111001110101101011000;
   assign mem[476543:476512] = 32'b00000010101000011010000011000000;
   assign mem[476575:476544] = 32'b00000100011011000111011000010000;
   assign mem[476607:476576] = 32'b11111001001110011001101011110000;
   assign mem[476639:476608] = 32'b00000010001000111111100001000100;
   assign mem[476671:476640] = 32'b11111001111101111110010100110000;
   assign mem[476703:476672] = 32'b11111100100010010111000000111100;
   assign mem[476735:476704] = 32'b00000001111100001001001011110010;
   assign mem[476767:476736] = 32'b11111010101000010000010101101000;
   assign mem[476799:476768] = 32'b00000101001101000101110000100000;
   assign mem[476831:476800] = 32'b00000100011001110001110001101000;
   assign mem[476863:476832] = 32'b00000010011001000000111001000100;
   assign mem[476895:476864] = 32'b00000101100111101101100100110000;
   assign mem[476927:476896] = 32'b00000011010111010000011011111000;
   assign mem[476959:476928] = 32'b11111100010001011000010001111100;
   assign mem[476991:476960] = 32'b11111100010111001011110000101100;
   assign mem[477023:476992] = 32'b00000001111110111100100010010010;
   assign mem[477055:477024] = 32'b00000101111110000011110001011000;
   assign mem[477087:477056] = 32'b00000001011111110111000000010110;
   assign mem[477119:477088] = 32'b11110000001001011110100011010000;
   assign mem[477151:477120] = 32'b00000101011111110000111111000000;
   assign mem[477183:477152] = 32'b11101111100001001110000100000000;
   assign mem[477215:477184] = 32'b00000001011011001110110000011100;
   assign mem[477247:477216] = 32'b00000100011011011001101100011000;
   assign mem[477279:477248] = 32'b11110001011010010100011101100000;
   assign mem[477311:477280] = 32'b00000011000001011100111101100000;
   assign mem[477343:477312] = 32'b00000011001100010111111111110100;
   assign mem[477375:477344] = 32'b11111000110010000110010010111000;
   assign mem[477407:477376] = 32'b00000100100111100000110111100000;
   assign mem[477439:477408] = 32'b11111100111100011110111111011100;
   assign mem[477471:477440] = 32'b11101010101101101010010001000000;
   assign mem[477503:477472] = 32'b11111110110000110100111101010000;
   assign mem[477535:477504] = 32'b11110111111000110111101111000000;
   assign mem[477567:477536] = 32'b11111011111111001001001110011000;
   assign mem[477599:477568] = 32'b00000111101010010101011000110000;
   assign mem[477631:477600] = 32'b11111100100010100011011111001000;
   assign mem[477663:477632] = 32'b11110010010100010010110111000000;
   assign mem[477695:477664] = 32'b00001101100110011011100010110000;
   assign mem[477727:477696] = 32'b11110111010001010100011100010000;
   assign mem[477759:477728] = 32'b00001000111101101111000110110000;
   assign mem[477791:477760] = 32'b00000011001011100010000100111100;
   assign mem[477823:477792] = 32'b00000001001010110011100001100100;
   assign mem[477855:477824] = 32'b00000011111001001000010110000000;
   assign mem[477887:477856] = 32'b00000001010101000101010111011110;
   assign mem[477919:477888] = 32'b11101110001010100000100001000000;
   assign mem[477951:477920] = 32'b00000010111001110101101110000100;
   assign mem[477983:477952] = 32'b11111111100110110100101001100011;
   assign mem[478015:477984] = 32'b11110100011110111101001010110000;
   assign mem[478047:478016] = 32'b00000011111000000010111011001000;
   assign mem[478079:478048] = 32'b11111110111101110010100100010000;
   assign mem[478111:478080] = 32'b00000001110100110010100011111100;
   assign mem[478143:478112] = 32'b11101101110000011001110101000000;
   assign mem[478175:478144] = 32'b11111111000010110001110111010000;
   assign mem[478207:478176] = 32'b00000101001010010010000101001000;
   assign mem[478239:478208] = 32'b11111001101001000111111101000000;
   assign mem[478271:478240] = 32'b00000010111001111101111111001000;
   assign mem[478303:478272] = 32'b00000001100011000010011000011110;
   assign mem[478335:478304] = 32'b11111010101010100100011011100000;
   assign mem[478367:478336] = 32'b00000101010100111101010011100000;
   assign mem[478399:478368] = 32'b11111100100110110101100010110000;
   assign mem[478431:478400] = 32'b11110001001000011111100011000000;
   assign mem[478463:478432] = 32'b00000000111111100100011111111101;
   assign mem[478495:478464] = 32'b00000010100111010001010101110100;
   assign mem[478527:478496] = 32'b11111100000011100010010010101100;
   assign mem[478559:478528] = 32'b00000001110010101011000110001100;
   assign mem[478591:478560] = 32'b11111000110101110111100001101000;
   assign mem[478623:478592] = 32'b11110111101101000001111000100000;
   assign mem[478655:478624] = 32'b00000011111100011011111110011000;
   assign mem[478687:478656] = 32'b11111110110110011001101111110010;
   assign mem[478719:478688] = 32'b00000011010000110001001011110100;
   assign mem[478751:478720] = 32'b11111011101101100111100010100000;
   assign mem[478783:478752] = 32'b11111111010111100100111000011011;
   assign mem[478815:478784] = 32'b00000101110001010010110101010000;
   assign mem[478847:478816] = 32'b00000000010010100101110000110001;
   assign mem[478879:478848] = 32'b00000010110000010000111100100000;
   assign mem[478911:478880] = 32'b11111100000010100101101100011000;
   assign mem[478943:478912] = 32'b11101111011100001110100100000000;
   assign mem[478975:478944] = 32'b11111101001011100010101011011000;
   assign mem[479007:478976] = 32'b11111110110000101001011101110000;
   assign mem[479039:479008] = 32'b00000001010010111101101101010100;
   assign mem[479071:479040] = 32'b11111100011011110000100111000000;
   assign mem[479103:479072] = 32'b00000010100000101101010010010100;
   assign mem[479135:479104] = 32'b11111000100010110100011101101000;
   assign mem[479167:479136] = 32'b11111111010000110000011111010001;
   assign mem[479199:479168] = 32'b00000000010000000001110100001101;
   assign mem[479231:479200] = 32'b00000001011001001111111001111000;
   assign mem[479263:479232] = 32'b11111110101000101011101111101000;
   assign mem[479295:479264] = 32'b00000000100111111101110111000111;
   assign mem[479327:479296] = 32'b11111111111101110010010011001101;
   assign mem[479359:479328] = 32'b00000010111111011011011101010100;
   assign mem[479391:479360] = 32'b11110110110111110000101101010000;
   assign mem[479423:479392] = 32'b11111111100000001110011101001111;
   assign mem[479455:479424] = 32'b11111000101101111101100010100000;
   assign mem[479487:479456] = 32'b11111101001110011100000001100100;
   assign mem[479519:479488] = 32'b00000011001101101110001110010100;
   assign mem[479551:479520] = 32'b11111000110110101111000000101000;
   assign mem[479583:479552] = 32'b11110101111011111000001110100000;
   assign mem[479615:479584] = 32'b00000000110110011110111110011110;
   assign mem[479647:479616] = 32'b00000010110101100000010001001100;
   assign mem[479679:479648] = 32'b00000100111000111111001001110000;
   assign mem[479711:479680] = 32'b00000111101111101101111111011000;
   assign mem[479743:479712] = 32'b00000010000101001110111110000000;
   assign mem[479775:479744] = 32'b11110110100101010110011000010000;
   assign mem[479807:479776] = 32'b11111110110000000001000010100000;
   assign mem[479839:479808] = 32'b11110101011000110000100001110000;
   assign mem[479871:479840] = 32'b00000000001000000111011100111010;
   assign mem[479903:479872] = 32'b00000111101010001110011000110000;
   assign mem[479935:479904] = 32'b00000011011010101100011000000000;
   assign mem[479967:479936] = 32'b11111010010001110111000001101000;
   assign mem[479999:479968] = 32'b00000011010001110010100000001100;
   assign mem[480031:480000] = 32'b00000101010010011000010100000000;
   assign mem[480063:480032] = 32'b00000011100111010100110110111100;
   assign mem[480095:480064] = 32'b00000011010010100101001011001000;
   assign mem[480127:480096] = 32'b11111110011110110111110110111110;
   assign mem[480159:480128] = 32'b11111000110000111111000100010000;
   assign mem[480191:480160] = 32'b00000000010010010111110010111101;
   assign mem[480223:480192] = 32'b00000100100100000011101100001000;
   assign mem[480255:480224] = 32'b11111011110100001011011000101000;
   assign mem[480287:480256] = 32'b00000011111101111001010001000100;
   assign mem[480319:480288] = 32'b11111101001001010100101001010000;
   assign mem[480351:480320] = 32'b00000101101001001100000111111000;
   assign mem[480383:480352] = 32'b11110110110011010111011001000000;
   assign mem[480415:480384] = 32'b00000101111010011011010101010000;
   assign mem[480447:480416] = 32'b00000010001010000100101110010000;
   assign mem[480479:480448] = 32'b11110110001100011111110001000000;
   assign mem[480511:480480] = 32'b11111111010100111101101011000000;
   assign mem[480543:480512] = 32'b00000100110000011011111010101000;
   assign mem[480575:480544] = 32'b11110000101010010110000110100000;
   assign mem[480607:480576] = 32'b00000001111110001110101011010100;
   assign mem[480639:480608] = 32'b11110110101101000001011001110000;
   assign mem[480671:480640] = 32'b11111010111100001110101101011000;
   assign mem[480703:480672] = 32'b00000001001101110101001001101000;
   assign mem[480735:480704] = 32'b11111001000111110101001100010000;
   assign mem[480767:480736] = 32'b11111100100000111011101100100100;
   assign mem[480799:480768] = 32'b00000101000100110100001100101000;
   assign mem[480831:480800] = 32'b11111111001101011001011001001011;
   assign mem[480863:480832] = 32'b11111100101100011101101100101100;
   assign mem[480895:480864] = 32'b00000001001100110000010110110100;
   assign mem[480927:480896] = 32'b00000000001110001111001011111001;
   assign mem[480959:480928] = 32'b00000101001111000000111001001000;
   assign mem[480991:480960] = 32'b00000100011101001100111011000000;
   assign mem[481023:480992] = 32'b00000001110111000011000110110100;
   assign mem[481055:481024] = 32'b00000011000001010010110010100100;
   assign mem[481087:481056] = 32'b00000001011001111100010010100000;
   assign mem[481119:481088] = 32'b11111100101111010000010011000100;
   assign mem[481151:481120] = 32'b11111100100101000000111011100100;
   assign mem[481183:481152] = 32'b11111110111101110011100101100010;
   assign mem[481215:481184] = 32'b00000001110011000100000111010000;
   assign mem[481247:481216] = 32'b11111110111010001110011111011100;
   assign mem[481279:481248] = 32'b11111101110101111010001001010100;
   assign mem[481311:481280] = 32'b00000111010000110101011011100000;
   assign mem[481343:481312] = 32'b11110011000001001010110000110000;
   assign mem[481375:481344] = 32'b00000010001111000001010000110100;
   assign mem[481407:481376] = 32'b00000110001010100011101111100000;
   assign mem[481439:481408] = 32'b11110100111011001010001001100000;
   assign mem[481471:481440] = 32'b00000101100101011111011010000000;
   assign mem[481503:481472] = 32'b11111100010110000011111001110100;
   assign mem[481535:481504] = 32'b11111011110100000000001101101000;
   assign mem[481567:481536] = 32'b11111010111011010101101101111000;
   assign mem[481599:481568] = 32'b11111110111001001001111001100100;
   assign mem[481631:481600] = 32'b11111101110101011111001100000000;
   assign mem[481663:481632] = 32'b11110101011110110011010101000000;
   assign mem[481695:481664] = 32'b11111100101011000101010010011000;
   assign mem[481727:481696] = 32'b00001000000111110000110000000000;
   assign mem[481759:481728] = 32'b00000000110001101101100111101001;
   assign mem[481791:481760] = 32'b11111110100100010001000100110110;
   assign mem[481823:481792] = 32'b00000100001111010100011001111000;
   assign mem[481855:481824] = 32'b00000110010000001111101000010000;
   assign mem[481887:481856] = 32'b11111101000100111000100110001000;
   assign mem[481919:481888] = 32'b11111100100100101001000000100000;
   assign mem[481951:481920] = 32'b00000001100000011100110010010000;
   assign mem[481983:481952] = 32'b00000010110101100110001000011100;
   assign mem[482015:481984] = 32'b00000100110100110001001000011000;
   assign mem[482047:482016] = 32'b11111111000010011111000110010100;
   assign mem[482079:482048] = 32'b11111110011011010010111101100100;
   assign mem[482111:482080] = 32'b11111011001000100011111111110000;
   assign mem[482143:482112] = 32'b00000010011001110110011011111100;
   assign mem[482175:482144] = 32'b11111010000011010000010010111000;
   assign mem[482207:482176] = 32'b00000001111110011100100010000000;
   assign mem[482239:482208] = 32'b11110111010011110111101010000000;
   assign mem[482271:482240] = 32'b00000100001011010110101100001000;
   assign mem[482303:482272] = 32'b00000001111101001001100100100000;
   assign mem[482335:482304] = 32'b11110110111001101000011001010000;
   assign mem[482367:482336] = 32'b00000111000110111001011110111000;
   assign mem[482399:482368] = 32'b11111111101101110110110010101011;
   assign mem[482431:482400] = 32'b00000011100100011110100100010000;
   assign mem[482463:482432] = 32'b00000001111000101010101110011110;
   assign mem[482495:482464] = 32'b11111110111100010100011001001000;
   assign mem[482527:482496] = 32'b00000100000101100000001000110000;
   assign mem[482559:482528] = 32'b00000001000000101100011110101010;
   assign mem[482591:482560] = 32'b00000100010101111101011011010000;
   assign mem[482623:482592] = 32'b00000110000001001110011010010000;
   assign mem[482655:482624] = 32'b00000110001100111100100001101000;
   assign mem[482687:482656] = 32'b00000001100110110100000010101000;
   assign mem[482719:482688] = 32'b11110010010110011100010100010000;
   assign mem[482751:482720] = 32'b00000001011110111101011101000110;
   assign mem[482783:482752] = 32'b00000010110001110011011001101000;
   assign mem[482815:482784] = 32'b11111100010101110100100101110000;
   assign mem[482847:482816] = 32'b00000011100010011000110101001000;
   assign mem[482879:482848] = 32'b11101111101000001100011001000000;
   assign mem[482911:482880] = 32'b11111000110000111001101101100000;
   assign mem[482943:482912] = 32'b00001011001101000101011001010000;
   assign mem[482975:482944] = 32'b00000110001100101101000100100000;
   assign mem[483007:482976] = 32'b11111111011110000001111110011110;
   assign mem[483039:483008] = 32'b00000101110110100101110111011000;
   assign mem[483071:483040] = 32'b11111101001011001110001010110000;
   assign mem[483103:483072] = 32'b11111111000001001000101001000001;
   assign mem[483135:483104] = 32'b00000000001110011110100111011001;
   assign mem[483167:483136] = 32'b00000001011011001101000111011010;
   assign mem[483199:483168] = 32'b11110011010010111001101011000000;
   assign mem[483231:483200] = 32'b00000001101101010011000010110010;
   assign mem[483263:483232] = 32'b00001001001100011011100100110000;
   assign mem[483295:483264] = 32'b00000011110101000100111101001000;
   assign mem[483327:483296] = 32'b11110110010001000000000110100000;
   assign mem[483359:483328] = 32'b00000000010100100100011011011111;
   assign mem[483391:483360] = 32'b11111000111011010001000000011000;
   assign mem[483423:483392] = 32'b00000101111110001100100010110000;
   assign mem[483455:483424] = 32'b11111010101100111001011101001000;
   assign mem[483487:483456] = 32'b00000010100111000110111101110100;
   assign mem[483519:483488] = 32'b00000001101001110111100100011100;
   assign mem[483551:483520] = 32'b00000011100101000111100010011100;
   assign mem[483583:483552] = 32'b00000100010010000011101110000000;
   assign mem[483615:483584] = 32'b00000010110100101001001111011100;
   assign mem[483647:483616] = 32'b00000111010001000100101011010000;
   assign mem[483679:483648] = 32'b11101101011000110110110011000000;
   assign mem[483711:483680] = 32'b11111110100101111110101011011110;
   assign mem[483743:483712] = 32'b00000101101000000000000001011000;
   assign mem[483775:483744] = 32'b11110011111001101000111100100000;
   assign mem[483807:483776] = 32'b00000000111110010010101111001111;
   assign mem[483839:483808] = 32'b11111000001011011001010001100000;
   assign mem[483871:483840] = 32'b11111100000111000111101001111100;
   assign mem[483903:483872] = 32'b00000001101010101011001100110100;
   assign mem[483935:483904] = 32'b00001001010111011101110010010000;
   assign mem[483967:483936] = 32'b00000001000010000101101011100010;
   assign mem[483999:483968] = 32'b11111111100111101111111000101000;
   assign mem[484031:484000] = 32'b11110101110101110100010100100000;
   assign mem[484063:484032] = 32'b00000011101011111100011100000100;
   assign mem[484095:484064] = 32'b00000000011001010001001101001010;
   assign mem[484127:484096] = 32'b11111001011011101000011110010000;
   assign mem[484159:484128] = 32'b11111101110111011101000001001000;
   assign mem[484191:484160] = 32'b00000011010110110001101111011000;
   assign mem[484223:484192] = 32'b00000000010000000101100100010011;
   assign mem[484255:484224] = 32'b00000001101001111000110100010110;
   assign mem[484287:484256] = 32'b00000000010111010100000001001111;
   assign mem[484319:484288] = 32'b11111101111000000011000101010000;
   assign mem[484351:484320] = 32'b11111111100011001110010101100100;
   assign mem[484383:484352] = 32'b00000100000100010000111111101000;
   assign mem[484415:484384] = 32'b11111011000010110110111011100000;
   assign mem[484447:484416] = 32'b11111010010100101110111111111000;
   assign mem[484479:484448] = 32'b11111011111111011010010100001000;
   assign mem[484511:484480] = 32'b00000010011101100010100101100000;
   assign mem[484543:484512] = 32'b00000011001100010011110010011000;
   assign mem[484575:484544] = 32'b00001000001001111011111011000000;
   assign mem[484607:484576] = 32'b11111001110111101111100011100000;
   assign mem[484639:484608] = 32'b11111100011111100001011101100100;
   assign mem[484671:484640] = 32'b11111010000011010111011010101000;
   assign mem[484703:484672] = 32'b00000111001001011111001111011000;
   assign mem[484735:484704] = 32'b00000001100010110000011000111010;
   assign mem[484767:484736] = 32'b11111100000010010111010001000100;
   assign mem[484799:484768] = 32'b11110111100101101110111001010000;
   assign mem[484831:484800] = 32'b11101101100000011101001001100000;
   assign mem[484863:484832] = 32'b11111111111110000010010000110111;
   assign mem[484895:484864] = 32'b11111111100011110110101011111110;
   assign mem[484927:484896] = 32'b00000011110111100011001100011000;
   assign mem[484959:484928] = 32'b11111010010011011010111010100000;
   assign mem[484991:484960] = 32'b00001001000010010110100111000000;
   assign mem[485023:484992] = 32'b11111100110110101010001000100000;
   assign mem[485055:485024] = 32'b11111011101010101111110101000000;
   assign mem[485087:485056] = 32'b00000110011001101010001000011000;
   assign mem[485119:485088] = 32'b11111100010001000001100011111000;
   assign mem[485151:485120] = 32'b11111111100100111110100011111010;
   assign mem[485183:485152] = 32'b00000110110100011100101010100000;
   assign mem[485215:485184] = 32'b00000110011001011011110110100000;
   assign mem[485247:485216] = 32'b11101110101011011011111011000000;
   assign mem[485279:485248] = 32'b11111111100101110001110011110111;
   assign mem[485311:485280] = 32'b11110110000000111001001011000000;
   assign mem[485343:485312] = 32'b00000011010101000000011111100000;
   assign mem[485375:485344] = 32'b00000100010010100000110110100000;
   assign mem[485407:485376] = 32'b11111110110000111111111011010010;
   assign mem[485439:485408] = 32'b11111110000101101011100010111110;
   assign mem[485471:485440] = 32'b11110100011011100111101011110000;
   assign mem[485503:485472] = 32'b00000001011110111000110010001110;
   assign mem[485535:485504] = 32'b00001001100110011100100110110000;
   assign mem[485567:485536] = 32'b00001010010101010110101110010000;
   assign mem[485599:485568] = 32'b11111000011000110100010100000000;
   assign mem[485631:485600] = 32'b00001010011001101011000010110000;
   assign mem[485663:485632] = 32'b11111010111000111010110010110000;
   assign mem[485695:485664] = 32'b11110101011101111101011001110000;
   assign mem[485727:485696] = 32'b00000011101000010111000011100000;
   assign mem[485759:485728] = 32'b11101001110101101101111011000000;
   assign mem[485791:485760] = 32'b11101101111000100110110100100000;
   assign mem[485823:485792] = 32'b00010000011010110111110010000000;
   assign mem[485855:485824] = 32'b00000000010000001000010000001010;
   assign mem[485887:485856] = 32'b00000101110110100111000110011000;
   assign mem[485919:485888] = 32'b00000110001100100001110101001000;
   assign mem[485951:485920] = 32'b11110100001000000000111111000000;
   assign mem[485983:485952] = 32'b11111001110010000000100010110000;
   assign mem[486015:485984] = 32'b00000101101110010011011000000000;
   assign mem[486047:486016] = 32'b11110011110001110000011011110000;
   assign mem[486079:486048] = 32'b00000111011110010010110100101000;
   assign mem[486111:486080] = 32'b00000010011101100000010011000000;
   assign mem[486143:486112] = 32'b11111110011111011101110001011100;
   assign mem[486175:486144] = 32'b11111100000011011111101001101100;
   assign mem[486207:486176] = 32'b11111101001001110011110101100100;
   assign mem[486239:486208] = 32'b11111110011100111000111000000100;
   assign mem[486271:486240] = 32'b00000010011101000110000111100000;
   assign mem[486303:486272] = 32'b11111110010101000001110010001100;
   assign mem[486335:486304] = 32'b11111111100011000001101111010110;
   assign mem[486367:486336] = 32'b00000000011110001100101101010111;
   assign mem[486399:486368] = 32'b00000010000100000110000010101000;
   assign mem[486431:486400] = 32'b00000001110010000001111010000100;
   assign mem[486463:486432] = 32'b00000110011111100001000000111000;
   assign mem[486495:486464] = 32'b00000101100010010111100001110000;
   assign mem[486527:486496] = 32'b00000100110001000111001110110000;
   assign mem[486559:486528] = 32'b11111101101100010000011011110100;
   assign mem[486591:486560] = 32'b00000100100110100011010100001000;
   assign mem[486623:486592] = 32'b00000011111100000100100000000100;
   assign mem[486655:486624] = 32'b11111110000001110110001111010010;
   assign mem[486687:486656] = 32'b11111100111001010011111111001100;
   assign mem[486719:486688] = 32'b11111010010010010111001000000000;
   assign mem[486751:486720] = 32'b00000101010000011000110110011000;
   assign mem[486783:486752] = 32'b11111010000100010011100110011000;
   assign mem[486815:486784] = 32'b11111110101100001111110000000010;
   assign mem[486847:486816] = 32'b00000111111110100111111001110000;
   assign mem[486879:486848] = 32'b11110100001110011100000110010000;
   assign mem[486911:486880] = 32'b11111110010011111011010000110010;
   assign mem[486943:486912] = 32'b00001000110000100001101010000000;
   assign mem[486975:486944] = 32'b00000100100010001001110100000000;
   assign mem[487007:486976] = 32'b00000001011000111010100110010010;
   assign mem[487039:487008] = 32'b11111010010100011001111111010000;
   assign mem[487071:487040] = 32'b11111101010100101111110000000100;
   assign mem[487103:487072] = 32'b11111001101001001010001000110000;
   assign mem[487135:487104] = 32'b11111111100001000101000110111101;
   assign mem[487167:487136] = 32'b00000111100010000111000110111000;
   assign mem[487199:487168] = 32'b11110011100000100100000010100000;
   assign mem[487231:487200] = 32'b00000110111011011101000000101000;
   assign mem[487263:487232] = 32'b00000011100100100000000110110000;
   assign mem[487295:487264] = 32'b11110110111010101000101001110000;
   assign mem[487327:487296] = 32'b00000110101100111011111111000000;
   assign mem[487359:487328] = 32'b11111110100010000001010111101000;
   assign mem[487391:487360] = 32'b11110001110010000011001001000000;
   assign mem[487423:487392] = 32'b00000111111111110011011100101000;
   assign mem[487455:487424] = 32'b00000101111111010000000011010000;
   assign mem[487487:487456] = 32'b00000000110111111111101011001101;
   assign mem[487519:487488] = 32'b00000101100010010001100010000000;
   assign mem[487551:487520] = 32'b11110110111001000111001110110000;
   assign mem[487583:487552] = 32'b11110110110010011111100000010000;
   assign mem[487615:487584] = 32'b00001000001011011011001011010000;
   assign mem[487647:487616] = 32'b11110101011110100110010111110000;
   assign mem[487679:487648] = 32'b00001000100001010001110010100000;
   assign mem[487711:487680] = 32'b00000010100011100100111010110000;
   assign mem[487743:487712] = 32'b00000011101111110110111101010100;
   assign mem[487775:487744] = 32'b00000011111110100010011111001000;
   assign mem[487807:487776] = 32'b11111110110010110110111000001110;
   assign mem[487839:487808] = 32'b00000001000000011100010101001010;
   assign mem[487871:487840] = 32'b11111110001001111011010001100110;
   assign mem[487903:487872] = 32'b00000011001011011111100100000100;
   assign mem[487935:487904] = 32'b11110011111011101001101011100000;
   assign mem[487967:487936] = 32'b00000000110110110001000111100011;
   assign mem[487999:487968] = 32'b11111110000111011111010000100110;
   assign mem[488031:488000] = 32'b00000101000000100110110000010000;
   assign mem[488063:488032] = 32'b00000011000101011011110011000000;
   assign mem[488095:488064] = 32'b00000100111011111010001110110000;
   assign mem[488127:488096] = 32'b11111111000111010000010100011111;
   assign mem[488159:488128] = 32'b11111010011001010001101010100000;
   assign mem[488191:488160] = 32'b11111110101010101110100001100110;
   assign mem[488223:488192] = 32'b00000110000000000011111000010000;
   assign mem[488255:488224] = 32'b11110011000011111001100110010000;
   assign mem[488287:488256] = 32'b00000001011111111010111011011000;
   assign mem[488319:488288] = 32'b11111111110100101101110100011001;
   assign mem[488351:488320] = 32'b00000011010011101001111000001100;
   assign mem[488383:488352] = 32'b00000010010100111110110011011100;
   assign mem[488415:488384] = 32'b00000000110010111000011100101010;
   assign mem[488447:488416] = 32'b11111111110110001010000110000010;
   assign mem[488479:488448] = 32'b11111001000101101110000011101000;
   assign mem[488511:488480] = 32'b00000001101100011101110011110100;
   assign mem[488543:488512] = 32'b00000000111111010110001100011101;
   assign mem[488575:488544] = 32'b11110011111100000011110000100000;
   assign mem[488607:488576] = 32'b00000001101100000011000011101100;
   assign mem[488639:488608] = 32'b11111111110000111000110011001111;
   assign mem[488671:488640] = 32'b00000010111101000001011011001100;
   assign mem[488703:488672] = 32'b11110011111110110110101000100000;
   assign mem[488735:488704] = 32'b11110101000001111111011011000000;
   assign mem[488767:488736] = 32'b00000101010000000110010011111000;
   assign mem[488799:488768] = 32'b11111011110010010111101011011000;
   assign mem[488831:488800] = 32'b00001000110100011011001000000000;
   assign mem[488863:488832] = 32'b00000001000101001101101101101000;
   assign mem[488895:488864] = 32'b11111111001111000111110010101110;
   assign mem[488927:488896] = 32'b00000101100110000011000110101000;
   assign mem[488959:488928] = 32'b11111110111001010101001101101100;
   assign mem[488991:488960] = 32'b11110101110100010010000111000000;
   assign mem[489023:488992] = 32'b00000000001100101101011110011101;
   assign mem[489055:489024] = 32'b11111001000000010100010100101000;
   assign mem[489087:489056] = 32'b00000110010110111010110000000000;
   assign mem[489119:489088] = 32'b11110111111011010000000111100000;
   assign mem[489151:489120] = 32'b00001000101100000010100110010000;
   assign mem[489183:489152] = 32'b00000100100101101100001010100000;
   assign mem[489215:489184] = 32'b11111001110001010000001111101000;
   assign mem[489247:489216] = 32'b00000110000101000111111000111000;
   assign mem[489279:489248] = 32'b11110111001111000001001101000000;
   assign mem[489311:489280] = 32'b11111110000111110010011010000010;
   assign mem[489343:489312] = 32'b11111011111111111100110001000000;
   assign mem[489375:489344] = 32'b00000011100110010000000010111100;
   assign mem[489407:489376] = 32'b00000010100011110001111000011100;
   assign mem[489439:489408] = 32'b11111101111001001100110100110100;
   assign mem[489471:489440] = 32'b11111111111010101000011101001001;
   assign mem[489503:489472] = 32'b00000001010111110011011111101000;
   assign mem[489535:489504] = 32'b11111010100000000010101000100000;
   assign mem[489567:489536] = 32'b11111000110111010110011000000000;
   assign mem[489599:489568] = 32'b11111010001011010011011110011000;
   assign mem[489631:489600] = 32'b11111111101100011001010110100110;
   assign mem[489663:489632] = 32'b11111010000111100111100011010000;
   assign mem[489695:489664] = 32'b00000000010010010101010010100011;
   assign mem[489727:489696] = 32'b00001000110000110000110011100000;
   assign mem[489759:489728] = 32'b11110001000000011010010010110000;
   assign mem[489791:489760] = 32'b00000110011111110100100001101000;
   assign mem[489823:489792] = 32'b11111110000011101001001001101100;
   assign mem[489855:489824] = 32'b11110000000001101111011110010000;
   assign mem[489887:489856] = 32'b00000010010111000010110100100100;
   assign mem[489919:489888] = 32'b11111000010000001100011011101000;
   assign mem[489951:489920] = 32'b11110110111011101111101100110000;
   assign mem[489983:489952] = 32'b00000000110100011011111001011110;
   assign mem[490015:489984] = 32'b00000011100101011111100011100100;
   assign mem[490047:490016] = 32'b00000011110100000101010100110000;
   assign mem[490079:490048] = 32'b11110111011100001010001010000000;
   assign mem[490111:490080] = 32'b00000110011100100101110001000000;
   assign mem[490143:490112] = 32'b00000011100010001111001100010000;
   assign mem[490175:490144] = 32'b11110000101010110000010110000000;
   assign mem[490207:490176] = 32'b00001000101010000010101001100000;
   assign mem[490239:490208] = 32'b11110111011011110010101010110000;
   assign mem[490271:490240] = 32'b00000100101001011100100101110000;
   assign mem[490303:490272] = 32'b00000011110100101110101001111100;
   assign mem[490335:490304] = 32'b00000111011010010111010011101000;
   assign mem[490367:490336] = 32'b00001001111010011011010101000000;
   assign mem[490399:490368] = 32'b11101100000100011001010100000000;
   assign mem[490431:490400] = 32'b00000101100100101101101001101000;
   assign mem[490463:490432] = 32'b00000010110101110011110101101100;
   assign mem[490495:490464] = 32'b11111011110001101100101111111000;
   assign mem[490527:490496] = 32'b00000010110001000110100111101100;
   assign mem[490559:490528] = 32'b11110001111001110100001010110000;
   assign mem[490591:490560] = 32'b00000110001001110101100010000000;
   assign mem[490623:490592] = 32'b11110011010001100101000101110000;
   assign mem[490655:490624] = 32'b11111100000000011100010100111000;
   assign mem[490687:490656] = 32'b00000101000011101011001110000000;
   assign mem[490719:490688] = 32'b11110110100101101001111100110000;
   assign mem[490751:490720] = 32'b00000010101110111010111101010000;
   assign mem[490783:490752] = 32'b11111111110001000010010100101100;
   assign mem[490815:490784] = 32'b00001110011111101010011110000000;
   assign mem[490847:490816] = 32'b11111011101100001111001100101000;
   assign mem[490879:490848] = 32'b11111011011101100111101100100000;
   assign mem[490911:490880] = 32'b11110000011111010000000110110000;
   assign mem[490943:490912] = 32'b00000100101000011001000000111000;
   assign mem[490975:490944] = 32'b11110111101111100111111100110000;
   assign mem[491007:490976] = 32'b11111001101101110001001011010000;
   assign mem[491039:491008] = 32'b00000100000001011101110110110000;
   assign mem[491071:491040] = 32'b11110101001011010011111111110000;
   assign mem[491103:491072] = 32'b11101101111110011010100001000000;
   assign mem[491135:491104] = 32'b00001001000011000100010010010000;
   assign mem[491167:491136] = 32'b11101101010000011101110000000000;
   assign mem[491199:491168] = 32'b00001000000100011011111101010000;
   assign mem[491231:491200] = 32'b00000000110001110100111100111100;
   assign mem[491263:491232] = 32'b11110110110001101011110101110000;
   assign mem[491295:491264] = 32'b11110110110000101110101110110000;
   assign mem[491327:491296] = 32'b00001000000010001001100011110000;
   assign mem[491359:491328] = 32'b11111110011011011110110001001000;
   assign mem[491391:491360] = 32'b11111110100011101100010001011010;
   assign mem[491423:491392] = 32'b11111101101101000110100101000000;
   assign mem[491455:491424] = 32'b11111110110100110110111111001010;
   assign mem[491487:491456] = 32'b11111110011111000001011011100010;
   assign mem[491519:491488] = 32'b11111110111101010100011100010000;
   assign mem[491551:491520] = 32'b00001000001001010101101011110000;
   assign mem[491583:491552] = 32'b11111011011001101101110001011000;
   assign mem[491615:491584] = 32'b00000101001000110001010000110000;
   assign mem[491647:491616] = 32'b11111010010111000010010101001000;
   assign mem[491679:491648] = 32'b11101111111011111111101101100000;
   assign mem[491711:491680] = 32'b00000101110100111101110011000000;
   assign mem[491743:491712] = 32'b11111110100111010010000111101100;
   assign mem[491775:491744] = 32'b00000010111111111101111101100100;
   assign mem[491807:491776] = 32'b00000001011111100110010000100000;
   assign mem[491839:491808] = 32'b11111111101111110010011000111010;
   assign mem[491871:491840] = 32'b11101001100001011011011001000000;
   assign mem[491903:491872] = 32'b00000110111110110100011111110000;
   assign mem[491935:491904] = 32'b00000100010111100111001100101000;
   assign mem[491967:491936] = 32'b00000010000010000101001000000000;
   assign mem[491999:491968] = 32'b11111011110100110110101001000000;
   assign mem[492031:492000] = 32'b11111110011110110011010010010000;
   assign mem[492063:492032] = 32'b11111010101100110101001000000000;
   assign mem[492095:492064] = 32'b11111010001100110011111000111000;
   assign mem[492127:492096] = 32'b00000011111101100001011000111000;
   assign mem[492159:492128] = 32'b00000000110001001011111011000100;
   assign mem[492191:492160] = 32'b11101111001101111110110001100000;
   assign mem[492223:492192] = 32'b00001001000010111011011001110000;
   assign mem[492255:492224] = 32'b00001100000010010101111110010000;
   assign mem[492287:492256] = 32'b11111011110111001001000110100000;
   assign mem[492319:492288] = 32'b00000100110011010100011000001000;
   assign mem[492351:492320] = 32'b11110101001010111001000001110000;
   assign mem[492383:492352] = 32'b11111101001000101011001000110000;
   assign mem[492415:492384] = 32'b11110011001101111000100110110000;
   assign mem[492447:492416] = 32'b11111110000110101011101000001100;
   assign mem[492479:492448] = 32'b00000000001000000100010110001110;
   assign mem[492511:492480] = 32'b00000001101000001101010100001110;
   assign mem[492543:492512] = 32'b00000110101011011111100100111000;
   assign mem[492575:492544] = 32'b00000111000100000001011010000000;
   assign mem[492607:492576] = 32'b11110110010110011000010010110000;
   assign mem[492639:492608] = 32'b00000101000111001101000100010000;
   assign mem[492671:492640] = 32'b11111000001110000011000101010000;
   assign mem[492703:492672] = 32'b00000100011101111011011000100000;
   assign mem[492735:492704] = 32'b00000001111010010000011101001010;
   assign mem[492767:492736] = 32'b11110011000110111110101001110000;
   assign mem[492799:492768] = 32'b11110110010010000000000111010000;
   assign mem[492831:492800] = 32'b00000011111100110111011110010100;
   assign mem[492863:492832] = 32'b11111111101000001001101110011000;
   assign mem[492895:492864] = 32'b00000001110100011111111110100000;
   assign mem[492927:492896] = 32'b11111011100101000111000011110000;
   assign mem[492959:492928] = 32'b00000010101110001001111011110100;
   assign mem[492991:492960] = 32'b11111011011010011001101111011000;
   assign mem[493023:492992] = 32'b00000011101100111001111111000100;
   assign mem[493055:493024] = 32'b11111111000100101000010011100111;
   assign mem[493087:493056] = 32'b11111101110001110111101101010000;
   assign mem[493119:493088] = 32'b11110111010010001010110100010000;
   assign mem[493151:493120] = 32'b00000011110111000100100111010000;
   assign mem[493183:493152] = 32'b11110110111000000101001001100000;
   assign mem[493215:493184] = 32'b11110110111101111010001011100000;
   assign mem[493247:493216] = 32'b00000110000101110101001010000000;
   assign mem[493279:493248] = 32'b11111100100100010010110010011000;
   assign mem[493311:493280] = 32'b00000110000010111010001000011000;
   assign mem[493343:493312] = 32'b11110111111010100001100001000000;
   assign mem[493375:493344] = 32'b11111101110101000110100101101000;
   assign mem[493407:493376] = 32'b00000110000010010001010011001000;
   assign mem[493439:493408] = 32'b11111011110001010010101010100000;
   assign mem[493471:493440] = 32'b00000000100010001011010011100101;
   assign mem[493503:493472] = 32'b11111101110111001100011001010100;
   assign mem[493535:493504] = 32'b11111110001111000000011001101010;
   assign mem[493567:493536] = 32'b00000001000110011011101101011010;
   assign mem[493599:493568] = 32'b11111110101101110000101100111000;
   assign mem[493631:493600] = 32'b11111111101000111001010111010100;
   assign mem[493663:493632] = 32'b00000000100010110000101010111000;
   assign mem[493695:493664] = 32'b11111111100100011010101101000011;
   assign mem[493727:493696] = 32'b11111110101101011010000010011010;
   assign mem[493759:493728] = 32'b11111011011111010101100001011000;
   assign mem[493791:493760] = 32'b00000111001011000000110101001000;
   assign mem[493823:493792] = 32'b11111001011111100001000011100000;
   assign mem[493855:493824] = 32'b11111001101101011111001011011000;
   assign mem[493887:493856] = 32'b00000010000000110100001011000100;
   assign mem[493919:493888] = 32'b11110011100001010100100101100000;
   assign mem[493951:493920] = 32'b00000000011100000010111011000001;
   assign mem[493983:493952] = 32'b00000000001101010010110000011101;
   assign mem[494015:493984] = 32'b11111110001000110101010000111110;
   assign mem[494047:494016] = 32'b11111111111100101000100011010100;
   assign mem[494079:494048] = 32'b11111100001011100100100100000000;
   assign mem[494111:494080] = 32'b11111111110100000000000000111111;
   assign mem[494143:494112] = 32'b00000111000001111100110001101000;
   assign mem[494175:494144] = 32'b00010011001100111111011100000000;
   assign mem[494207:494176] = 32'b11110001111001001110001010000000;
   assign mem[494239:494208] = 32'b00001000110000011101100001010000;
   assign mem[494271:494240] = 32'b11111000101001100100110000101000;
   assign mem[494303:494272] = 32'b11101100110110100110001111100000;
   assign mem[494335:494304] = 32'b11110011000100011101111000000000;
   assign mem[494367:494336] = 32'b11110100101110100101010011010000;
   assign mem[494399:494368] = 32'b00000110011111001010001111000000;
   assign mem[494431:494400] = 32'b00001000001110001010100100100000;
   assign mem[494463:494432] = 32'b11110001001110111100110011100000;
   assign mem[494495:494464] = 32'b11111000000011010010111000100000;
   assign mem[494527:494496] = 32'b00001000000000100010110111100000;
   assign mem[494559:494528] = 32'b11111011100001100010100101110000;
   assign mem[494591:494560] = 32'b11111111111110011100111101111000;
   assign mem[494623:494592] = 32'b00000110000110111101111111000000;
   assign mem[494655:494624] = 32'b11111100010011100101110001100000;
   assign mem[494687:494656] = 32'b00000000000110111010101000001011;
   assign mem[494719:494688] = 32'b11111011101100101001011000000000;
   assign mem[494751:494720] = 32'b00000001100011101111100100000100;
   assign mem[494783:494752] = 32'b00000011101100101010100000010100;
   assign mem[494815:494784] = 32'b00001010111100010111101000000000;
   assign mem[494847:494816] = 32'b11111000000010110111111000100000;
   assign mem[494879:494848] = 32'b00000010011011011000110010011100;
   assign mem[494911:494880] = 32'b11111011010111101000000111000000;
   assign mem[494943:494912] = 32'b11111011011110000001110110000000;
   assign mem[494975:494944] = 32'b11110101100001010110101111100000;
   assign mem[495007:494976] = 32'b11111110011101100101110110111100;
   assign mem[495039:495008] = 32'b00000001011110110111110111001110;
   assign mem[495071:495040] = 32'b11110110000000101011111001010000;
   assign mem[495103:495072] = 32'b00000110110010111010101101001000;
   assign mem[495135:495104] = 32'b00001101011101010011110001010000;
   assign mem[495167:495136] = 32'b11110000110111100010001001100000;
   assign mem[495199:495168] = 32'b00001000100001101110000001010000;
   assign mem[495231:495200] = 32'b11111011110011100000011011010000;
   assign mem[495263:495232] = 32'b11111100100001000010011111011000;
   assign mem[495295:495264] = 32'b11111010111010000011000001101000;
   assign mem[495327:495296] = 32'b11110111101101100101101100010000;
   assign mem[495359:495328] = 32'b00000110001011010010110111101000;
   assign mem[495391:495360] = 32'b11110011000001011010100001010000;
   assign mem[495423:495392] = 32'b11111000000111110010000010110000;
   assign mem[495455:495424] = 32'b00011011000010001001100101100000;
   assign mem[495487:495456] = 32'b11110111010101100111111010010000;
   assign mem[495519:495488] = 32'b00000100101011010001101001010000;
   assign mem[495551:495520] = 32'b11110100000011110110110000100000;
   assign mem[495583:495552] = 32'b00000000101100001001010011111110;
   assign mem[495615:495584] = 32'b11110101101111100001111100010000;
   assign mem[495647:495616] = 32'b11110010110000010111100001000000;
   assign mem[495679:495648] = 32'b00000110111110011001101011111000;
   assign mem[495711:495680] = 32'b11101000101101000010111010000000;
   assign mem[495743:495712] = 32'b00000010111001101011110100110000;
   assign mem[495775:495744] = 32'b00010100100101100100100011100000;
   assign mem[495807:495776] = 32'b11111000001101110011101010100000;
   assign mem[495839:495808] = 32'b00001010110100001011111101010000;
   assign mem[495871:495840] = 32'b11110100101111111100000011000000;
   assign mem[495903:495872] = 32'b11110100010000100110001011110000;
   assign mem[495935:495904] = 32'b11110100110000000010111010110000;
   assign mem[495967:495936] = 32'b11110110110111001011100000110000;
   assign mem[495999:495968] = 32'b11111111110001101000111010001011;
   assign mem[496031:496000] = 32'b11111000011110000011000101101000;
   assign mem[496063:496032] = 32'b00000101111101000101111010101000;
   assign mem[496095:496064] = 32'b00001111011111011000010010010000;
   assign mem[496127:496096] = 32'b11111100101011111100101010101000;
   assign mem[496159:496128] = 32'b00000100001110011100010100100000;
   assign mem[496191:496160] = 32'b11111001111000111001111000110000;
   assign mem[496223:496192] = 32'b11111101100111011111011111010000;
   assign mem[496255:496224] = 32'b11111011001001001001111100110000;
   assign mem[496287:496256] = 32'b11110101111111101100101011110000;
   assign mem[496319:496288] = 32'b00000001000001000011010010011100;
   assign mem[496351:496320] = 32'b11111111110100011011111000010001;
   assign mem[496383:496352] = 32'b11111010000001001001110010011000;
   assign mem[496415:496384] = 32'b11110000000011101101001110100000;
   assign mem[496447:496416] = 32'b00000110100000001101100000100000;
   assign mem[496479:496448] = 32'b11111100001110101100001100001100;
   assign mem[496511:496480] = 32'b11111111111111101100000000000111;
   assign mem[496543:496512] = 32'b11111011111001101000111110100000;
   assign mem[496575:496544] = 32'b11111001001100111000101111111000;
   assign mem[496607:496576] = 32'b00001000100010000001110010100000;
   assign mem[496639:496608] = 32'b11111001110111011010110010111000;
   assign mem[496671:496640] = 32'b00000001100011010011100111110100;
   assign mem[496703:496672] = 32'b00000011110011111101110011110000;
   assign mem[496735:496704] = 32'b00001000110111111110111010100000;
   assign mem[496767:496736] = 32'b11111010000111111111010001111000;
   assign mem[496799:496768] = 32'b00000110010111111001010000011000;
   assign mem[496831:496800] = 32'b11111100111000001101010101011000;
   assign mem[496863:496832] = 32'b00000011110110000100010111000100;
   assign mem[496895:496864] = 32'b11110010101011111011100010110000;
   assign mem[496927:496896] = 32'b00000000001000001110000111000001;
   assign mem[496959:496928] = 32'b11110110011000101101101101010000;
   assign mem[496991:496960] = 32'b11111111010110001001000011000001;
   assign mem[497023:496992] = 32'b11111110101110101100111001001010;
   assign mem[497055:497024] = 32'b00000011000011111100010111100100;
   assign mem[497087:497056] = 32'b11110110110100010111011101110000;
   assign mem[497119:497088] = 32'b00001101011110110100000101110000;
   assign mem[497151:497120] = 32'b11111000111111000010111111100000;
   assign mem[497183:497152] = 32'b11111110101101100101011000100100;
   assign mem[497215:497184] = 32'b11110000001110111111111110100000;
   assign mem[497247:497216] = 32'b00000011001010110101110101101000;
   assign mem[497279:497248] = 32'b00000110011000001011000110110000;
   assign mem[497311:497280] = 32'b00001000111000101000001011100000;
   assign mem[497343:497312] = 32'b00000000010101111011100010010010;
   assign mem[497375:497344] = 32'b00000111010011111100000111101000;
   assign mem[497407:497376] = 32'b11111011100101110101011010011000;
   assign mem[497439:497408] = 32'b00000001101100101111010010101100;
   assign mem[497471:497440] = 32'b11110010100100011101001110010000;
   assign mem[497503:497472] = 32'b00000001010111001010101101001100;
   assign mem[497535:497504] = 32'b00000010101001111000101111011000;
   assign mem[497567:497536] = 32'b11111111111110001001000001000110;
   assign mem[497599:497568] = 32'b11111000101010111000011110110000;
   assign mem[497631:497600] = 32'b00001111011011000101010101000000;
   assign mem[497663:497632] = 32'b11111111101000111100000011001100;
   assign mem[497695:497664] = 32'b11111101111101000111101011110000;
   assign mem[497727:497696] = 32'b00000101111010010010000110001000;
   assign mem[497759:497728] = 32'b11111101101101000001001010000100;
   assign mem[497791:497760] = 32'b11111111010011110011000111000000;
   assign mem[497823:497792] = 32'b00000100000000001001111110100000;
   assign mem[497855:497824] = 32'b11110111100011010011010110000000;
   assign mem[497887:497856] = 32'b00000010010011111011010000101100;
   assign mem[497919:497888] = 32'b11101100110011001100101000100000;
   assign mem[497951:497920] = 32'b11101110111100110011000111100000;
   assign mem[497983:497952] = 32'b11111110110011110111000110101010;
   assign mem[498015:497984] = 32'b00000000110000100001101100000000;
   assign mem[498047:498016] = 32'b11111101100111101000000100011000;
   assign mem[498079:498048] = 32'b00001101100110110100010101110000;
   assign mem[498111:498080] = 32'b00000000011000001000001000001100;
   assign mem[498143:498112] = 32'b11101101001001110000110100000000;
   assign mem[498175:498144] = 32'b11111010001110100010111000100000;
   assign mem[498207:498176] = 32'b00000010100010110010101111101100;
   assign mem[498239:498208] = 32'b00001001000111101110101101100000;
   assign mem[498271:498240] = 32'b11111110000100101110110100111100;
   assign mem[498303:498272] = 32'b00000000010111111110001111111110;
   assign mem[498335:498304] = 32'b00001101000000100010010111010000;
   assign mem[498367:498336] = 32'b00000000000111100000011110010110;
   assign mem[498399:498368] = 32'b00000110000101111000100010100000;
   assign mem[498431:498400] = 32'b00000001111101100000001101101110;
   assign mem[498463:498432] = 32'b00000001000000001100100000110110;
   assign mem[498495:498464] = 32'b11110011001000110101010000000000;
   assign mem[498527:498496] = 32'b00000000101010000101010000000000;
   assign mem[498559:498528] = 32'b11110100110010110000000000010000;
   assign mem[498591:498560] = 32'b00000100110000011000001111111000;
   assign mem[498623:498592] = 32'b11111000011100100010010100011000;
   assign mem[498655:498624] = 32'b11110101010110011000010010010000;
   assign mem[498687:498656] = 32'b00000101111000100011110011101000;
   assign mem[498719:498688] = 32'b11110010101001110000010110000000;
   assign mem[498751:498720] = 32'b00000011010001000100101000101000;
   assign mem[498783:498752] = 32'b00000010011000111010110010111000;
   assign mem[498815:498784] = 32'b11111100011010100010110101100000;
   assign mem[498847:498816] = 32'b00000011110100101010110001111100;
   assign mem[498879:498848] = 32'b11111011101101100100000111011000;
   assign mem[498911:498880] = 32'b11110010111100110111010110000000;
   assign mem[498943:498912] = 32'b00001000110111010110000100000000;
   assign mem[498975:498944] = 32'b00000000011011110101110100010011;
   assign mem[499007:498976] = 32'b11111101001001111100111011111000;
   assign mem[499039:499008] = 32'b00000010101011001011011101010100;
   assign mem[499071:499040] = 32'b11111011110001111001011100010000;
   assign mem[499103:499072] = 32'b11110011001010001110011000000000;
   assign mem[499135:499104] = 32'b11111100000111110000100110110100;
   assign mem[499167:499136] = 32'b11111111111101010101011010110001;
   assign mem[499199:499168] = 32'b00001001011101011100000001000000;
   assign mem[499231:499200] = 32'b11101110110001111011110100000000;
   assign mem[499263:499232] = 32'b11111100110111011100110001111000;
   assign mem[499295:499264] = 32'b00000010001110101001010100011100;
   assign mem[499327:499296] = 32'b00000000111101011000101100000001;
   assign mem[499359:499328] = 32'b00000001100100111110000010111010;
   assign mem[499391:499360] = 32'b11111011011111111010001101001000;
   assign mem[499423:499392] = 32'b11111010011001011011110100111000;
   assign mem[499455:499424] = 32'b11111000000000111110101001001000;
   assign mem[499487:499456] = 32'b00000001010011010010011100101010;
   assign mem[499519:499488] = 32'b00001001100101100010100010000000;
   assign mem[499551:499520] = 32'b11111110011000011000111111111010;
   assign mem[499583:499552] = 32'b11111110011101100101100000000010;
   assign mem[499615:499584] = 32'b11111101010011101000111100110100;
   assign mem[499647:499616] = 32'b00000100000010000101100110001000;
   assign mem[499679:499648] = 32'b00000010100111010101011011001000;
   assign mem[499711:499680] = 32'b11111111001100101000100000011000;
   assign mem[499743:499712] = 32'b11111111101011110110000011110110;
   assign mem[499775:499744] = 32'b00000000001011100011011101101000;
   assign mem[499807:499776] = 32'b11111111001100100100101110000000;
   assign mem[499839:499808] = 32'b11111101001110111110000000001100;
   assign mem[499871:499840] = 32'b11111010100010011001001100001000;
   assign mem[499903:499872] = 32'b11111011111101111111010111011000;
   assign mem[499935:499904] = 32'b00000001011110110001110010011110;
   assign mem[499967:499936] = 32'b11111110111111101100001011001100;
   assign mem[499999:499968] = 32'b00000010101000000010011000111000;
   assign mem[500031:500000] = 32'b11111010011100110010100000011000;
   assign mem[500063:500032] = 32'b11111010011000001000111111010000;
   assign mem[500095:500064] = 32'b00000101111001000001011100000000;
   assign mem[500127:500096] = 32'b11111101111111010101100000010100;
   assign mem[500159:500128] = 32'b00000011100101000101001111100000;
   assign mem[500191:500160] = 32'b00001011101110110000101001000000;
   assign mem[500223:500192] = 32'b11101100000111111000100111100000;
   assign mem[500255:500224] = 32'b11110101100111101100011110100000;
   assign mem[500287:500256] = 32'b00000110111101011110111100010000;
   assign mem[500319:500288] = 32'b00000001000111101011000011000000;
   assign mem[500351:500320] = 32'b00000010001111011111010110100100;
   assign mem[500383:500352] = 32'b00001000101001110011110101110000;
   assign mem[500415:500384] = 32'b00000111011101010001011001101000;
   assign mem[500447:500416] = 32'b11111110100110101110010101001100;
   assign mem[500479:500448] = 32'b11111100011111011101001011100100;
   assign mem[500511:500480] = 32'b11111000011000011010111100000000;
   assign mem[500543:500512] = 32'b00000000000000001110010000111011;
   assign mem[500575:500544] = 32'b00001001110000110010010010010000;
   assign mem[500607:500576] = 32'b11111011101100100010100100001000;
   assign mem[500639:500608] = 32'b00000000111111001001000011011001;
   assign mem[500671:500640] = 32'b11111110000110101110100000111010;
   assign mem[500703:500672] = 32'b00000101010001110100011010101000;
   assign mem[500735:500704] = 32'b11111000101100011011011110101000;
   assign mem[500767:500736] = 32'b00000101101101010001111000101000;
   assign mem[500799:500768] = 32'b11111101010011010111000101011000;
   assign mem[500831:500800] = 32'b00000010010110001001001111100100;
   assign mem[500863:500832] = 32'b00000111101101100110110101011000;
   assign mem[500895:500864] = 32'b00010101101000110110101100100000;
   assign mem[500927:500896] = 32'b11101110101111101101010010100000;
   assign mem[500959:500928] = 32'b00000010010101111011001111101100;
   assign mem[500991:500960] = 32'b11111111000001011110000111000010;
   assign mem[501023:500992] = 32'b11110011111010000000110100100000;
   assign mem[501055:501024] = 32'b11101111100011101000100011000000;
   assign mem[501087:501056] = 32'b11111000011011111011010111101000;
   assign mem[501119:501088] = 32'b11111000001001001110000001010000;
   assign mem[501151:501120] = 32'b11110101011100000100101111100000;
   assign mem[501183:501152] = 32'b11111011110111010000000000101000;
   assign mem[501215:501184] = 32'b11101110100100111111000110100000;
   assign mem[501247:501216] = 32'b00000011110111111010110111010100;
   assign mem[501279:501248] = 32'b11111111111011111001010110010111;
   assign mem[501311:501280] = 32'b11111111011011110110010001001110;
   assign mem[501343:501312] = 32'b11111111110100111101001001010100;
   assign mem[501375:501344] = 32'b00000011101011010010001000101100;
   assign mem[501407:501376] = 32'b00000011000000101100110001100000;
   assign mem[501439:501408] = 32'b00000000010111100011100000111100;
   assign mem[501471:501440] = 32'b00000000100101010011110011100010;
   assign mem[501503:501472] = 32'b00000101101000101111011110010000;
   assign mem[501535:501504] = 32'b00000110111100110111010101010000;
   assign mem[501567:501536] = 32'b11111010000001101101100011110000;
   assign mem[501599:501568] = 32'b00000111101001000101001010000000;
   assign mem[501631:501600] = 32'b11110110010011100010000101010000;
   assign mem[501663:501632] = 32'b11111101000000000101001001100000;
   assign mem[501695:501664] = 32'b00000001111000010000111010000000;
   assign mem[501727:501696] = 32'b00000001001101101000010110001000;
   assign mem[501759:501728] = 32'b11110100010011011001011000110000;
   assign mem[501791:501760] = 32'b00000111011001100000011100010000;
   assign mem[501823:501792] = 32'b11110001011111101111011100110000;
   assign mem[501855:501824] = 32'b11110101111110010111011111100000;
   assign mem[501887:501856] = 32'b00000110101101011001001000110000;
   assign mem[501919:501888] = 32'b11101110111101000111110110000000;
   assign mem[501951:501920] = 32'b00000111110000101101101000011000;
   assign mem[501983:501952] = 32'b00000011101110010011001011010000;
   assign mem[502015:501984] = 32'b11111011000101110100111011001000;
   assign mem[502047:502016] = 32'b00000100100111101010100011011000;
   assign mem[502079:502048] = 32'b11110111010111011010111111110000;
   assign mem[502111:502080] = 32'b00000000010110110100011111100100;
   assign mem[502143:502112] = 32'b11111100101011000100101100001100;
   assign mem[502175:502144] = 32'b11110011101011000010011010110000;
   assign mem[502207:502176] = 32'b00000100110000001111000111011000;
   assign mem[502239:502208] = 32'b11111011110111001100100101010000;
   assign mem[502271:502240] = 32'b00000100000010101001000110001000;
   assign mem[502303:502272] = 32'b11111100011110101011101111000100;
   assign mem[502335:502304] = 32'b11111100010101101101110000110100;
   assign mem[502367:502336] = 32'b11111111010111010110010100010100;
   assign mem[502399:502368] = 32'b00000011101111110100000100101100;
   assign mem[502431:502400] = 32'b11111111010111001011001100101000;
   assign mem[502463:502432] = 32'b00000111110111001011010011101000;
   assign mem[502495:502464] = 32'b00000110011000101100000011111000;
   assign mem[502527:502496] = 32'b11111010001101110101101111011000;
   assign mem[502559:502528] = 32'b11111111100111111011100010000001;
   assign mem[502591:502560] = 32'b11110110111000101010001010100000;
   assign mem[502623:502592] = 32'b00000000000001000101100110101101;
   assign mem[502655:502624] = 32'b11111100011111100110010000101000;
   assign mem[502687:502656] = 32'b11111100011011100110101001110000;
   assign mem[502719:502688] = 32'b11111101010010000100100111110000;
   assign mem[502751:502720] = 32'b00000011011001101001100000001000;
   assign mem[502783:502752] = 32'b11111011100011011001111101011000;
   assign mem[502815:502784] = 32'b11111010011011110001000010110000;
   assign mem[502847:502816] = 32'b00000001000100111110100100000000;
   assign mem[502879:502848] = 32'b11111101100011001010001010001100;
   assign mem[502911:502880] = 32'b00000010101101001111011000011100;
   assign mem[502943:502912] = 32'b00000010010101001001000010010000;
   assign mem[502975:502944] = 32'b11111111001000011001110101001010;
   assign mem[503007:502976] = 32'b00000000110001011101101110111100;
   assign mem[503039:503008] = 32'b11111100111101011111100111010100;
   assign mem[503071:503040] = 32'b00000010100111011001101000010100;
   assign mem[503103:503072] = 32'b00001100000111011101110010100000;
   assign mem[503135:503104] = 32'b00010100000110000010011101000000;
   assign mem[503167:503136] = 32'b11110110000110110110001100000000;
   assign mem[503199:503168] = 32'b00000000111001100110101100110110;
   assign mem[503231:503200] = 32'b11110000111101110011001000100000;
   assign mem[503263:503232] = 32'b11111010110000101010110000001000;
   assign mem[503295:503264] = 32'b11111011111011110000001010101000;
   assign mem[503327:503296] = 32'b11111001100111000111011100110000;
   assign mem[503359:503328] = 32'b11111100010011111000011001001100;
   assign mem[503391:503360] = 32'b11110001000110100011010111000000;
   assign mem[503423:503392] = 32'b00001001000101100110010001100000;
   assign mem[503455:503424] = 32'b00001010000101110101001000100000;
   assign mem[503487:503456] = 32'b11110110101100101101100100010000;
   assign mem[503519:503488] = 32'b00000101010111110110110010011000;
   assign mem[503551:503520] = 32'b11110110111100110011111110110000;
   assign mem[503583:503552] = 32'b11111001001001000010111010010000;
   assign mem[503615:503584] = 32'b11110101111010100001111010010000;
   assign mem[503647:503616] = 32'b11111100001111111000000001011100;
   assign mem[503679:503648] = 32'b00000000110100011001011000110010;
   assign mem[503711:503680] = 32'b11110011100001101010110101100000;
   assign mem[503743:503712] = 32'b00001101011111111101111011100000;
   assign mem[503775:503744] = 32'b00001110010011000111100100010000;
   assign mem[503807:503776] = 32'b11111010111110001001100100001000;
   assign mem[503839:503808] = 32'b00001000110010000111011110000000;
   assign mem[503871:503840] = 32'b11111001000010110010001001011000;
   assign mem[503903:503872] = 32'b11111001000111100000101010000000;
   assign mem[503935:503904] = 32'b11111101110110101110111110001000;
   assign mem[503967:503936] = 32'b11110111110100101010001111110000;
   assign mem[503999:503968] = 32'b00000011111010001011110011101000;
   assign mem[504031:504000] = 32'b00000110101111100100110101110000;
   assign mem[504063:504032] = 32'b00001000001000110001110000100000;
   assign mem[504095:504064] = 32'b00000101001111110110111000010000;
   assign mem[504127:504096] = 32'b11111000011000000000001111100000;
   assign mem[504159:504128] = 32'b00000000010010000011110001100010;
   assign mem[504191:504160] = 32'b11111000100011101110000011111000;
   assign mem[504223:504192] = 32'b00001001010001000000111001110000;
   assign mem[504255:504224] = 32'b11111010101111100000011100110000;
   assign mem[504287:504256] = 32'b11111111000100100110100110101010;
   assign mem[504319:504288] = 32'b11110111111110110101000010000000;
   assign mem[504351:504320] = 32'b11111111111001100100011100100000;
   assign mem[504383:504352] = 32'b00000010000010000001011100100100;
   assign mem[504415:504384] = 32'b00000111011001000101000001101000;
   assign mem[504447:504416] = 32'b11111100110111010011111101011100;
   assign mem[504479:504448] = 32'b00000011100011101001101110001000;
   assign mem[504511:504480] = 32'b11110110001011101101111100010000;
   assign mem[504543:504512] = 32'b00000000001001011001101101101100;
   assign mem[504575:504544] = 32'b11110101101011111101001111010000;
   assign mem[504607:504576] = 32'b11111000101101001000000110101000;
   assign mem[504639:504608] = 32'b00000011000101111111001010111100;
   assign mem[504671:504640] = 32'b00000011001110101000000110000000;
   assign mem[504703:504672] = 32'b00000101000010100111110011100000;
   assign mem[504735:504704] = 32'b00000100010101101100110100111000;
   assign mem[504767:504736] = 32'b11111100000001000101111101000100;
   assign mem[504799:504768] = 32'b00000011011011111110001111101100;
   assign mem[504831:504800] = 32'b11111101111111001110101101110100;
   assign mem[504863:504832] = 32'b11111010111011101000001011110000;
   assign mem[504895:504864] = 32'b11111111011010001010011011111001;
   assign mem[504927:504896] = 32'b11111101111001011101101011111000;
   assign mem[504959:504928] = 32'b11111111110100101110110110010100;
   assign mem[504991:504960] = 32'b11110111000011001110101111010000;
   assign mem[505023:504992] = 32'b00001001011011111111100100110000;
   assign mem[505055:505024] = 32'b00001110111100100101101011110000;
   assign mem[505087:505056] = 32'b11110011000010111000100111110000;
   assign mem[505119:505088] = 32'b00001010101101010010100001110000;
   assign mem[505151:505120] = 32'b11110111011011100010111111110000;
   assign mem[505183:505152] = 32'b11111100101011011110101101100100;
   assign mem[505215:505184] = 32'b11111011110010001101011111000000;
   assign mem[505247:505216] = 32'b11110110010111111101110011110000;
   assign mem[505279:505248] = 32'b11111111111000110010001101000000;
   assign mem[505311:505280] = 32'b11110101111111000001111010010000;
   assign mem[505343:505312] = 32'b00000100000000000001100111010000;
   assign mem[505375:505344] = 32'b11111100011111000111001111000100;
   assign mem[505407:505376] = 32'b00000011011011001010101001001100;
   assign mem[505439:505408] = 32'b00000000000000101000011101011100;
   assign mem[505471:505440] = 32'b00000000011000010111010000100100;
   assign mem[505503:505472] = 32'b00000011010000011001101000101000;
   assign mem[505535:505504] = 32'b11110111100100001001001010000000;
   assign mem[505567:505536] = 32'b00000101100000110111101111100000;
   assign mem[505599:505568] = 32'b11111100111011000100110101111100;
   assign mem[505631:505600] = 32'b11111100111111101100011011000100;
   assign mem[505663:505632] = 32'b00000011101010100011111011101100;
   assign mem[505695:505664] = 32'b00000010100010001101101111001100;
   assign mem[505727:505696] = 32'b11110100101010111101101101000000;
   assign mem[505759:505728] = 32'b00000110111000110111001100000000;
   assign mem[505791:505760] = 32'b11111000011010100000010000101000;
   assign mem[505823:505792] = 32'b11110001111111000001111110100000;
   assign mem[505855:505824] = 32'b00000100010000111011111000010000;
   assign mem[505887:505856] = 32'b11111111100111000100010110011010;
   assign mem[505919:505888] = 32'b00001011110000010010010001000000;
   assign mem[505951:505920] = 32'b11101100011100101110111000100000;
   assign mem[505983:505952] = 32'b00001001010101010100000011010000;
   assign mem[506015:505984] = 32'b00000001101001010101010011011100;
   assign mem[506047:506016] = 32'b00000111001001100001101100110000;
   assign mem[506079:506048] = 32'b11111011110111000111000110001000;
   assign mem[506111:506080] = 32'b11111001001110110010011001100000;
   assign mem[506143:506112] = 32'b00000010011111011101011101001100;
   assign mem[506175:506144] = 32'b11110010010110101011101000010000;
   assign mem[506207:506176] = 32'b00001000111011000000110010110000;
   assign mem[506239:506208] = 32'b11110111000110101000001110110000;
   assign mem[506271:506240] = 32'b11111101011010100110010111001000;
   assign mem[506303:506272] = 32'b00000111001110101100110111110000;
   assign mem[506335:506304] = 32'b00001000101100101001111110110000;
   assign mem[506367:506336] = 32'b11110100001101010101011100100000;
   assign mem[506399:506368] = 32'b00000100010001100110010010011000;
   assign mem[506431:506400] = 32'b00000000011101110000011011101110;
   assign mem[506463:506432] = 32'b11111000001101010110000101100000;
   assign mem[506495:506464] = 32'b11111000001111001011000000011000;
   assign mem[506527:506496] = 32'b11110100110100000101111110010000;
   assign mem[506559:506528] = 32'b00000001101101000100101110010110;
   assign mem[506591:506560] = 32'b00000010110011011110111010100000;
   assign mem[506623:506592] = 32'b11111111100111000001000000011101;
   assign mem[506655:506624] = 32'b11111100111011101000110000011000;
   assign mem[506687:506656] = 32'b11111111101000111001101000101011;
   assign mem[506719:506688] = 32'b11111101110001011011100001000000;
   assign mem[506751:506720] = 32'b00000010011110010100011101110000;
   assign mem[506783:506752] = 32'b00000010110111010111001111000000;
   assign mem[506815:506784] = 32'b00000010110111010111000011010100;
   assign mem[506847:506816] = 32'b11111110011100101101011000011100;
   assign mem[506879:506848] = 32'b00000000011000111010101111101110;
   assign mem[506911:506880] = 32'b00000011101010000011100101101100;
   assign mem[506943:506912] = 32'b00000000110101000110010110011011;
   assign mem[506975:506944] = 32'b00000111101110101011111111111000;
   assign mem[507007:506976] = 32'b00000010001001110111110111010100;
   assign mem[507039:507008] = 32'b00000000101001111010110110110101;
   assign mem[507071:507040] = 32'b11111001001000101001111101101000;
   assign mem[507103:507072] = 32'b11111110101100001101111101111000;
   assign mem[507135:507104] = 32'b00000011000101001011101101000000;
   assign mem[507167:507136] = 32'b11111110111001001010010101101010;
   assign mem[507199:507168] = 32'b11111101111101010101000110010100;
   assign mem[507231:507200] = 32'b00000110001101110010100100000000;
   assign mem[507263:507232] = 32'b11111011010101001101110110100000;
   assign mem[507295:507264] = 32'b00000011111000000000000000101100;
   assign mem[507327:507296] = 32'b00000001000001100010001100110110;
   assign mem[507359:507328] = 32'b11111111010111011011011001110101;
   assign mem[507391:507360] = 32'b00000011010100011010110010111100;
   assign mem[507423:507392] = 32'b11110101001101101011100101110000;
   assign mem[507455:507424] = 32'b11101111101000001011001001100000;
   assign mem[507487:507456] = 32'b00000011101101010110111111111000;
   assign mem[507519:507488] = 32'b11111011000100101000111000100000;
   assign mem[507551:507520] = 32'b11111100101100001101001101101100;
   assign mem[507583:507552] = 32'b11101011010001000001010010100000;
   assign mem[507615:507584] = 32'b11111100111011100000000011110000;
   assign mem[507647:507616] = 32'b00001001010100010010101110010000;
   assign mem[507679:507648] = 32'b11111000100001010101001011010000;
   assign mem[507711:507680] = 32'b00001000010110000100001110110000;
   assign mem[507743:507712] = 32'b00000111101110011010000010011000;
   assign mem[507775:507744] = 32'b11110100011111100100111111110000;
   assign mem[507807:507776] = 32'b00000100010101001001111011100000;
   assign mem[507839:507808] = 32'b11110111101010110111010001100000;
   assign mem[507871:507840] = 32'b11110110001100101110111001010000;
   assign mem[507903:507872] = 32'b00000011111101111000111111010100;
   assign mem[507935:507904] = 32'b00000100010010000110010010100000;
   assign mem[507967:507936] = 32'b11110000110011100111110010010000;
   assign mem[507999:507968] = 32'b11111111011011101000010001001101;
   assign mem[508031:508000] = 32'b00001011100010010100111110000000;
   assign mem[508063:508032] = 32'b11101010101000101100101000000000;
   assign mem[508095:508064] = 32'b11111000100010101100001110111000;
   assign mem[508127:508096] = 32'b11111100000010110010000100011100;
   assign mem[508159:508128] = 32'b00001011101010101001110101110000;
   assign mem[508191:508160] = 32'b11111110010111010100111110111000;
   assign mem[508223:508192] = 32'b00001010101110000001001110000000;
   assign mem[508255:508224] = 32'b00000111000111110000001111101000;
   assign mem[508287:508256] = 32'b11110110000001101010000111010000;
   assign mem[508319:508288] = 32'b00000110011001010000100011100000;
   assign mem[508351:508320] = 32'b11111011001111110011001010110000;
   assign mem[508383:508352] = 32'b00000000000110100111001001000100;
   assign mem[508415:508384] = 32'b11111000010001111100111011100000;
   assign mem[508447:508416] = 32'b00000011100010100001010110101100;
   assign mem[508479:508448] = 32'b00000000101110010110001101111111;
   assign mem[508511:508480] = 32'b00000011011110110010011011111000;
   assign mem[508543:508512] = 32'b00000010011110111010001111010000;
   assign mem[508575:508544] = 32'b00001001000000001011110000100000;
   assign mem[508607:508576] = 32'b11111001110101101010110111100000;
   assign mem[508639:508608] = 32'b00001000010000001110100011100000;
   assign mem[508671:508640] = 32'b11110110110001100010011110010000;
   assign mem[508703:508672] = 32'b00000011010011111101011101010000;
   assign mem[508735:508704] = 32'b11111100011110100100011101000100;
   assign mem[508767:508736] = 32'b00000101100001011000101001000000;
   assign mem[508799:508768] = 32'b11111011001110000101001100110000;
   assign mem[508831:508800] = 32'b00000011010011011011101101000000;
   assign mem[508863:508832] = 32'b00000001011001100000000010011100;
   assign mem[508895:508864] = 32'b00000010001000101111110111010000;
   assign mem[508927:508896] = 32'b11111110010111110111010111100010;
   assign mem[508959:508928] = 32'b11110111110001010101011100110000;
   assign mem[508991:508960] = 32'b11111010101111010001100010011000;
   assign mem[509023:508992] = 32'b11111010001110100000000110100000;
   assign mem[509055:509024] = 32'b11111000010111100101101100101000;
   assign mem[509087:509056] = 32'b00001001111101011000100101010000;
   assign mem[509119:509088] = 32'b11111001101100111100111100011000;
   assign mem[509151:509120] = 32'b11111111011111111001101111111001;
   assign mem[509183:509152] = 32'b11111010110001010111000110011000;
   assign mem[509215:509184] = 32'b11111100111111110011100101001000;
   assign mem[509247:509216] = 32'b00000011000100111100001011111000;
   assign mem[509279:509248] = 32'b11110111101001111001110101110000;
   assign mem[509311:509280] = 32'b00000001011110011101101011110000;
   assign mem[509343:509312] = 32'b00000000110010011001110010010011;
   assign mem[509375:509344] = 32'b11111011100000110111001011110000;
   assign mem[509407:509376] = 32'b00000100111010011100100101011000;
   assign mem[509439:509408] = 32'b11111110001101111001000011110100;
   assign mem[509471:509440] = 32'b11111111011101110001101111000011;
   assign mem[509503:509472] = 32'b00000100000100111100101001001000;
   assign mem[509535:509504] = 32'b11111101001101010010100111111100;
   assign mem[509567:509536] = 32'b11111100101110000011101001101000;
   assign mem[509599:509568] = 32'b11111010101010100101110001100000;
   assign mem[509631:509600] = 32'b00000010011010010001100100010000;
   assign mem[509663:509632] = 32'b00000001011101001000001011000100;
   assign mem[509695:509664] = 32'b11111000000010001000101010000000;
   assign mem[509727:509696] = 32'b00000100101001011100010101101000;
   assign mem[509759:509728] = 32'b11111111000111011011011011000110;
   assign mem[509791:509760] = 32'b11111010110011101011010100010000;
   assign mem[509823:509792] = 32'b00000011001010001101001001110000;
   assign mem[509855:509824] = 32'b00001000100010111011110101000000;
   assign mem[509887:509856] = 32'b11111100000111010011010100100000;
   assign mem[509919:509888] = 32'b00000111100110000110100110100000;
   assign mem[509951:509920] = 32'b11111011110001011001110011000000;
   assign mem[509983:509952] = 32'b11111101111000110000011010111100;
   assign mem[510015:509984] = 32'b11110111110001110010111011010000;
   assign mem[510047:510016] = 32'b11110100101000001101100010000000;
   assign mem[510079:510048] = 32'b11111100101000110111101001001100;
   assign mem[510111:510080] = 32'b11101111001100010100111111000000;
   assign mem[510143:510112] = 32'b00000110000010111011110000001000;
   assign mem[510175:510144] = 32'b00000110001100011101110110111000;
   assign mem[510207:510176] = 32'b00000010010111001000011011110000;
   assign mem[510239:510208] = 32'b11111011010111101100010101001000;
   assign mem[510271:510240] = 32'b11111000001100000110110110000000;
   assign mem[510303:510272] = 32'b11111111001100110111010000011010;
   assign mem[510335:510304] = 32'b11101110111111011100101011000000;
   assign mem[510367:510336] = 32'b00000111001101001001100010001000;
   assign mem[510399:510368] = 32'b00000000110101000111111011100111;
   assign mem[510431:510400] = 32'b11110100110100001001001010010000;
   assign mem[510463:510432] = 32'b11111111110101011001110111111111;
   assign mem[510495:510464] = 32'b00000011110111000011110100001000;
   assign mem[510527:510496] = 32'b00000101101010000010011100011000;
   assign mem[510559:510528] = 32'b11111110100101111101001011110000;
   assign mem[510591:510560] = 32'b00000010100011001110010011100100;
   assign mem[510623:510592] = 32'b00000000010011000100111011011011;
   assign mem[510655:510624] = 32'b11110001110111101101100010000000;
   assign mem[510687:510656] = 32'b00001010101000100101101000100000;
   assign mem[510719:510688] = 32'b11111111011100100110110010010010;
   assign mem[510751:510720] = 32'b00001010100011011010110101010000;
   assign mem[510783:510752] = 32'b11111011111000100100111000111000;
   assign mem[510815:510784] = 32'b00001010001100001000100010110000;
   assign mem[510847:510816] = 32'b11110010001101011010101000010000;
   assign mem[510879:510848] = 32'b00001010100101100110011111010000;
   assign mem[510911:510880] = 32'b11111110101110111110100011110100;
   assign mem[510943:510912] = 32'b00000001111110110001001110111010;
   assign mem[510975:510944] = 32'b11110101111101011111110000010000;
   assign mem[511007:510976] = 32'b11110110111000000000110001000000;
   assign mem[511039:511008] = 32'b11111001000011010000111111000000;
   assign mem[511071:511040] = 32'b00000100101111010101110111111000;
   assign mem[511103:511072] = 32'b11111101100101011010110001100100;
   assign mem[511135:511104] = 32'b00000101010111101110100101101000;
   assign mem[511167:511136] = 32'b00000101001010011100101010000000;
   assign mem[511199:511168] = 32'b11111101010111111010000110000000;
   assign mem[511231:511200] = 32'b00000010110100011001111000101000;
   assign mem[511263:511232] = 32'b11110101110101111101100111010000;
   assign mem[511295:511264] = 32'b11110110110101011110000111110000;
   assign mem[511327:511296] = 32'b11111100010111101111101100010000;
   assign mem[511359:511328] = 32'b11111111110001011000101110101101;
   assign mem[511391:511360] = 32'b11110011111011010000010110000000;
   assign mem[511423:511392] = 32'b00000001110001001101001111001000;
   assign mem[511455:511424] = 32'b11111111100010010001101111100110;
   assign mem[511487:511456] = 32'b11111011101111010100100000000000;
   assign mem[511519:511488] = 32'b00001001001010100011000011000000;
   assign mem[511551:511520] = 32'b00000011011110110001011010110100;
   assign mem[511583:511552] = 32'b11101111010101011110100101100000;
   assign mem[511615:511584] = 32'b11111000010101000011010010000000;
   assign mem[511647:511616] = 32'b11111101110010111000111101000000;
   assign mem[511679:511648] = 32'b00001011101000000101000101110000;
   assign mem[511711:511680] = 32'b11111000010101000010000000000000;
   assign mem[511743:511712] = 32'b11111110110100101100110111111000;
   assign mem[511775:511744] = 32'b11110011000110100110001011000000;
   assign mem[511807:511776] = 32'b11111101001011111010110000001100;
   assign mem[511839:511808] = 32'b11111101110110111111111000010000;
   assign mem[511871:511840] = 32'b00001000000110011000001100010000;
   assign mem[511903:511872] = 32'b11110111101111000100001000100000;
   assign mem[511935:511904] = 32'b11111001101011100100010100010000;
   assign mem[511967:511936] = 32'b00000010101010110010101110010000;
   assign mem[511999:511968] = 32'b11111111101011001100101101000010;


endmodule
